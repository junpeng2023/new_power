module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net962;
 wire net208;
 wire net966;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire clknet_0_clk;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net45;
 wire net289;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net963;
 wire net964;
 wire net965;
 wire net967;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net797;
 wire clknet_1_0__leaf_net797;
 wire clknet_1_1__leaf_net797;
 wire clknet_0_net796;
 wire clknet_1_0__leaf_net796;
 wire clknet_1_1__leaf_net796;
 wire clknet_0_net795;
 wire clknet_1_0__leaf_net795;
 wire clknet_1_1__leaf_net795;
 wire clknet_0_net777;
 wire clknet_1_0__leaf_net777;
 wire clknet_1_1__leaf_net777;
 wire clknet_0_net567;
 wire clknet_1_0__leaf_net567;
 wire clknet_1_1__leaf_net567;
 wire clknet_0_net590;
 wire clknet_1_0__leaf_net590;
 wire clknet_1_1__leaf_net590;
 wire clknet_0_net571;
 wire clknet_1_0__leaf_net571;
 wire clknet_1_1__leaf_net571;
 wire clknet_0_net568;
 wire clknet_1_0__leaf_net568;
 wire clknet_1_1__leaf_net568;
 wire clknet_0_net776;
 wire clknet_1_0__leaf_net776;
 wire clknet_1_1__leaf_net776;
 wire clknet_0_net775;
 wire clknet_1_0__leaf_net775;
 wire clknet_1_1__leaf_net775;
 wire clknet_0_net886;
 wire clknet_1_0__leaf_net886;
 wire clknet_1_1__leaf_net886;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net401;
 wire clknet_1_0__leaf_net401;
 wire clknet_1_1__leaf_net401;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net758;
 wire clknet_1_0__leaf_net758;
 wire clknet_1_1__leaf_net758;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net608;
 wire clknet_1_0__leaf_net608;
 wire clknet_1_1__leaf_net608;
 wire clknet_0_net493;
 wire clknet_1_0__leaf_net493;
 wire clknet_1_1__leaf_net493;
 wire clknet_0_net704;
 wire clknet_1_0__leaf_net704;
 wire clknet_1_1__leaf_net704;
 wire clknet_0_net508;
 wire clknet_1_0__leaf_net508;
 wire clknet_1_1__leaf_net508;
 wire clknet_0_net492;
 wire clknet_1_0__leaf_net492;
 wire clknet_1_1__leaf_net492;
 wire clknet_0_net488;
 wire clknet_1_0__leaf_net488;
 wire clknet_1_1__leaf_net488;
 wire clknet_0_net757;
 wire clknet_1_0__leaf_net757;
 wire clknet_1_1__leaf_net757;
 wire clknet_0_net739;
 wire clknet_1_0__leaf_net739;
 wire clknet_1_1__leaf_net739;
 wire clknet_0_net738;
 wire clknet_1_0__leaf_net738;
 wire clknet_1_1__leaf_net738;
 wire clknet_0_net266;
 wire clknet_1_0__leaf_net266;
 wire clknet_1_1__leaf_net266;
 wire clknet_0_net370;
 wire clknet_1_0__leaf_net370;
 wire clknet_1_1__leaf_net370;
 wire clknet_0_net881;
 wire clknet_1_0__leaf_net881;
 wire clknet_1_1__leaf_net881;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net707;
 wire clknet_1_0__leaf_net707;
 wire clknet_1_1__leaf_net707;
 wire clknet_0_net331;
 wire clknet_1_0__leaf_net331;
 wire clknet_1_1__leaf_net331;
 wire clknet_0_net706;
 wire clknet_1_0__leaf_net706;
 wire clknet_1_1__leaf_net706;
 wire clknet_0_net247;
 wire clknet_1_0__leaf_net247;
 wire clknet_1_1__leaf_net247;
 wire clknet_0_net217;
 wire clknet_1_0__leaf_net217;
 wire clknet_1_1__leaf_net217;
 wire clknet_0_net439;
 wire clknet_1_0__leaf_net439;
 wire clknet_1_1__leaf_net439;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net394;
 wire clknet_1_0__leaf_net394;
 wire clknet_1_1__leaf_net394;
 wire clknet_0_net329;
 wire clknet_1_0__leaf_net329;
 wire clknet_1_1__leaf_net329;
 wire clknet_0_net447;
 wire clknet_1_0__leaf_net447;
 wire clknet_1_1__leaf_net447;
 wire clknet_0_net432;
 wire clknet_1_0__leaf_net432;
 wire clknet_1_1__leaf_net432;
 wire clknet_0_net358;
 wire clknet_1_0__leaf_net358;
 wire clknet_1_1__leaf_net358;
 wire clknet_0_net344;
 wire clknet_1_0__leaf_net344;
 wire clknet_1_1__leaf_net344;
 wire clknet_0_net330;
 wire clknet_1_0__leaf_net330;
 wire clknet_1_1__leaf_net330;
 wire clknet_0_net240;
 wire clknet_1_0__leaf_net240;
 wire clknet_1_1__leaf_net240;
 wire clknet_0_net342;
 wire clknet_1_0__leaf_net342;
 wire clknet_1_1__leaf_net342;
 wire clknet_0_net241;
 wire clknet_1_0__leaf_net241;
 wire clknet_1_1__leaf_net241;
 wire clknet_0_net219;
 wire clknet_1_0__leaf_net219;
 wire clknet_1_1__leaf_net219;
 wire clknet_0_net256;
 wire clknet_1_0__leaf_net256;
 wire clknet_1_1__leaf_net256;
 wire clknet_0_net218;
 wire clknet_1_0__leaf_net218;
 wire clknet_1_1__leaf_net218;
 wire clknet_0_net234;
 wire clknet_1_0__leaf_net234;
 wire clknet_1_1__leaf_net234;
 wire clknet_0_net232;
 wire clknet_1_0__leaf_net232;
 wire clknet_1_1__leaf_net232;
 wire clknet_0_net454;
 wire clknet_1_0__leaf_net454;
 wire clknet_1_1__leaf_net454;
 wire clknet_0_net456;
 wire clknet_1_0__leaf_net456;
 wire clknet_1_1__leaf_net456;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net239;
 wire clknet_1_0__leaf_net239;
 wire clknet_1_1__leaf_net239;
 wire clknet_0_net254;
 wire clknet_1_0__leaf_net254;
 wire clknet_1_1__leaf_net254;
 wire net207;
 wire net209;
 wire net320;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net981;
 wire net982;
 wire net983;
 wire net1007;
 wire net1008;

 sky130_fd_sc_hd__or3b_2 c100 (.A(net10),
    .B(net30),
    .C_N(net29),
    .X(net36));
 sky130_fd_sc_hd__or2b_2 c101 (.A(net20),
    .B_N(net916),
    .X(net37));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net826),
    .A1(net30),
    .A2(net37),
    .A3(net26),
    .S0(net35),
    .S1(net25),
    .X(net38));
 sky130_fd_sc_hd__nand3_1 c103 (.A(net27),
    .B(net31),
    .C(net38),
    .Y(net39));
 sky130_fd_sc_hd__and3_1 c104 (.A(net30),
    .B(net20),
    .C(net35),
    .X(net40));
 sky130_fd_sc_hd__nor3_1 c105 (.A(net40),
    .B(net39),
    .C(net37),
    .Y(net41));
 sky130_fd_sc_hd__a211o_1 c106 (.A1(net41),
    .A2(net37),
    .B1(net36),
    .C1(net45),
    .X(net42));
 sky130_fd_sc_hd__a211oi_1 c107 (.A1(net33),
    .A2(net40),
    .B1(net35),
    .C1(net42),
    .Y(net43));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net39),
    .A1(net41),
    .A2(net29),
    .A3(net40),
    .S0(net30),
    .S1(net35),
    .X(net44));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net42),
    .A1(net44),
    .A2(net39),
    .A3(net37),
    .S0(net25),
    .X(net908));
 sky130_fd_sc_hd__inv_4 c110 (.A(net645),
    .Y(net46));
 sky130_fd_sc_hd__buf_1 c111 (.A(net645),
    .X(net47));
 sky130_fd_sc_hd__nand2_2 c112 (.A(net837),
    .B(net24),
    .Y(net898));
 sky130_fd_sc_hd__nand2b_1 c113 (.A_N(net857),
    .B(net18),
    .Y(net48));
 sky130_fd_sc_hd__and2_1 c114 (.A(net40),
    .B(net817),
    .X(net49));
 sky130_fd_sc_hd__buf_16 c115 (.A(net665),
    .X(net910));
 sky130_fd_sc_hd__and2b_1 c116 (.A_N(net840),
    .B(net32),
    .X(net50));
 sky130_fd_sc_hd__and2b_1 c117 (.A_N(net823),
    .B(net35),
    .X(net51));
 sky130_fd_sc_hd__nor3b_2 c118 (.A(net51),
    .B(net38),
    .C_N(net48),
    .Y(net52));
 sky130_fd_sc_hd__nand3b_1 c119 (.A_N(net38),
    .B(net898),
    .C(net52),
    .Y(net53));
 sky130_fd_sc_hd__inv_2 c120 (.A(net665),
    .Y(net54));
 sky130_fd_sc_hd__nand2b_2 c121 (.A_N(net52),
    .B(net49),
    .Y(net55));
 sky130_fd_sc_hd__or3b_2 c122 (.A(net46),
    .B(net50),
    .C_N(net40),
    .X(net925));
 sky130_fd_sc_hd__nand3_2 c123 (.A(net51),
    .B(net55),
    .C(net908),
    .Y(net56));
 sky130_fd_sc_hd__a221oi_1 c124 (.A1(net32),
    .A2(net55),
    .B1(net51),
    .B2(net24),
    .C1(net925),
    .Y(net57));
 sky130_fd_sc_hd__and3_1 c125 (.A(net50),
    .B(net51),
    .C(net52),
    .X(net888));
 sky130_fd_sc_hd__a221o_1 c126 (.A1(net55),
    .A2(net916),
    .B1(net898),
    .B2(net56),
    .C1(net692),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 c127 (.A(net708),
    .X(net59));
 sky130_fd_sc_hd__and3_1 c128 (.A(net59),
    .B(net46),
    .C(net692),
    .X(net60));
 sky130_fd_sc_hd__nand3b_4 c129 (.A_N(net48),
    .B(net52),
    .C(net60),
    .Y(net61));
 sky130_fd_sc_hd__a211o_1 c130 (.A1(net53),
    .A2(net60),
    .B1(net61),
    .C1(net18),
    .X(net906));
 sky130_fd_sc_hd__or3b_1 c131 (.A(net60),
    .B(net61),
    .C_N(net917),
    .X(net62));
 sky130_fd_sc_hd__nor2_2 c132 (.A(net821),
    .B(net815),
    .Y(net63));
 sky130_fd_sc_hd__and2b_2 c133 (.A_N(net869),
    .B(net815),
    .X(net64));
 sky130_fd_sc_hd__nand2_1 c134 (.A(net952),
    .B(net823),
    .Y(net65));
 sky130_fd_sc_hd__and2b_4 c135 (.A_N(net822),
    .B(net952),
    .X(net872));
 sky130_fd_sc_hd__or2b_4 c136 (.A(net65),
    .B_N(net872),
    .X(net66));
 sky130_fd_sc_hd__or3_1 c137 (.A(net812),
    .B(net868),
    .C(net952),
    .X(net67));
 sky130_fd_sc_hd__and2b_2 c138 (.A_N(net819),
    .B(net823),
    .X(net907));
 sky130_fd_sc_hd__and3_4 c139 (.A(net814),
    .B(net67),
    .C(net948),
    .X(net68));
 sky130_fd_sc_hd__and3_4 c140 (.A(net813),
    .B(net67),
    .C(net948),
    .X(net69));
 sky130_fd_sc_hd__a221oi_4 c141 (.A1(net68),
    .A2(net823),
    .B1(net832),
    .B2(net952),
    .C1(net949),
    .Y(net70));
 sky130_fd_sc_hd__nand2b_1 c142 (.A_N(net823),
    .B(net949),
    .Y(net71));
 sky130_fd_sc_hd__and2b_1 c143 (.A_N(net66),
    .B(net65),
    .X(net72));
 sky130_fd_sc_hd__nand2_2 c144 (.A(net65),
    .B(net68),
    .Y(net73));
 sky130_fd_sc_hd__a211oi_2 c145 (.A1(net870),
    .A2(net868),
    .B1(net948),
    .C1(net952),
    .Y(net74));
 sky130_fd_sc_hd__a211o_4 c146 (.A1(net854),
    .A2(net66),
    .B1(net868),
    .C1(net948),
    .X(net75));
 sky130_fd_sc_hd__or3_1 c147 (.A(net74),
    .B(net73),
    .C(net948),
    .X(net76));
 sky130_fd_sc_hd__and3_4 c148 (.A(net75),
    .B(net948),
    .C(net72),
    .X(net77));
 sky130_fd_sc_hd__mux4_2 c149 (.A0(net67),
    .A1(net77),
    .A2(net72),
    .A3(net872),
    .S0(net68),
    .S1(net813),
    .X(net78));
 sky130_fd_sc_hd__a221o_4 c150 (.A1(net78),
    .A2(net74),
    .B1(net76),
    .B2(net77),
    .C1(net948),
    .X(net79));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net77),
    .A1(net78),
    .A2(net952),
    .A3(net79),
    .S0(net948),
    .S1(net76),
    .X(net80));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net76),
    .A1(net66),
    .A2(net77),
    .A3(net939),
    .S0(net73),
    .S1(net79),
    .X(net81));
 sky130_fd_sc_hd__nand3_4 c153 (.A(net69),
    .B(net821),
    .C(net79),
    .Y(net82));
 sky130_fd_sc_hd__and2b_2 c154 (.A_N(net820),
    .B(net823),
    .X(net83));
 sky130_fd_sc_hd__nand2_2 c155 (.A(net816),
    .B(net79),
    .Y(net84));
 sky130_fd_sc_hd__or2b_2 c156 (.A(net846),
    .B_N(net70),
    .X(net85));
 sky130_fd_sc_hd__nor2_2 c157 (.A(net971),
    .B(net938),
    .Y(net904));
 sky130_fd_sc_hd__nor2_4 c158 (.A(net85),
    .B(net938),
    .Y(net927));
 sky130_fd_sc_hd__and2_1 c159 (.A(net937),
    .B(net872),
    .X(net86));
 sky130_fd_sc_hd__or3b_4 c160 (.A(net86),
    .B(net289),
    .C_N(net949),
    .X(net87));
 sky130_fd_sc_hd__a211oi_4 c161 (.A1(net837),
    .A2(net83),
    .B1(net827),
    .C1(net938),
    .Y(net88));
 sky130_fd_sc_hd__nor3_1 c162 (.A(net842),
    .B(net84),
    .C(net937),
    .Y(net89));
 sky130_fd_sc_hd__nand2_2 c163 (.A(net838),
    .B(net71),
    .Y(net90));
 sky130_fd_sc_hd__nor2b_1 c164 (.A(net839),
    .B_N(net79),
    .Y(net91));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net828),
    .A1(net89),
    .A2(net90),
    .A3(net86),
    .S0(net937),
    .S1(net838),
    .X(net92));
 sky130_fd_sc_hd__or3_1 c166 (.A(net89),
    .B(net834),
    .C(net937),
    .X(net93));
 sky130_fd_sc_hd__a221o_1 c167 (.A1(net71),
    .A2(net86),
    .B1(net938),
    .B2(net949),
    .C1(net937),
    .X(net94));
 sky130_fd_sc_hd__nand3b_4 c168 (.A_N(net73),
    .B(net91),
    .C(net939),
    .Y(net95));
 sky130_fd_sc_hd__nand2b_1 c169 (.A_N(net91),
    .B(net73),
    .Y(net96));
 sky130_fd_sc_hd__mux4_1 c170 (.A0(net831),
    .A1(net835),
    .A2(net96),
    .A3(net837),
    .S0(net937),
    .S1(net86),
    .X(net97));
 sky130_fd_sc_hd__or2_1 c171 (.A(net96),
    .B(net95),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net93),
    .A1(net96),
    .A2(net97),
    .A3(net937),
    .S0(net872),
    .S1(net971),
    .X(net99));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net99),
    .A1(net971),
    .A2(net98),
    .A3(net88),
    .S0(net73),
    .S1(net839),
    .X(net100));
 sky130_fd_sc_hd__a221o_4 c174 (.A1(net100),
    .A2(net839),
    .B1(net95),
    .B2(net938),
    .C1(net949),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net101),
    .A1(net99),
    .A2(net71),
    .A3(net97),
    .S0(net85),
    .S1(net100),
    .X(net883));
 sky130_fd_sc_hd__nand2b_1 c176 (.A_N(net865),
    .B(net840),
    .Y(net102));
 sky130_fd_sc_hd__buf_1 c177 (.A(net699),
    .X(net103));
 sky130_fd_sc_hd__nand2_2 c178 (.A(net827),
    .B(net953),
    .Y(net104));
 sky130_fd_sc_hd__nor3_1 c179 (.A(net102),
    .B(net953),
    .C(net69),
    .Y(net105));
 sky130_fd_sc_hd__and2_1 c180 (.A(net941),
    .B(net88),
    .X(net106));
 sky130_fd_sc_hd__and2_0 c181 (.A(net104),
    .B(net850),
    .X(net107));
 sky130_fd_sc_hd__nand3b_1 c182 (.A_N(net864),
    .B(net104),
    .C(net953),
    .Y(net108));
 sky130_fd_sc_hd__and2b_1 c183 (.A_N(net93),
    .B(net104),
    .X(net109));
 sky130_fd_sc_hd__nand3b_1 c184 (.A_N(net850),
    .B(net970),
    .C(net954),
    .Y(net110));
 sky130_fd_sc_hd__inv_1 c185 (.A(net699),
    .Y(net111));
 sky130_fd_sc_hd__a221o_2 c186 (.A1(net104),
    .A2(net853),
    .B1(net953),
    .B2(net110),
    .C1(net82),
    .X(net112));
 sky130_fd_sc_hd__a211o_1 c187 (.A1(net112),
    .A2(net105),
    .B1(net860),
    .C1(net953),
    .X(net113));
 sky130_fd_sc_hd__a221o_1 c188 (.A1(net111),
    .A2(net113),
    .B1(net864),
    .B2(net107),
    .C1(net953),
    .X(net114));
 sky130_fd_sc_hd__and3b_1 c189 (.A_N(net110),
    .B(net112),
    .C(net951),
    .X(net115));
 sky130_fd_sc_hd__a211oi_1 c190 (.A1(net840),
    .A2(net841),
    .B1(net112),
    .C1(net954),
    .Y(net116));
 sky130_fd_sc_hd__a221oi_2 c191 (.A1(net82),
    .A2(net116),
    .B1(net108),
    .B2(net112),
    .C1(net953),
    .Y(net117));
 sky130_fd_sc_hd__a221oi_4 c192 (.A1(net113),
    .A2(net104),
    .B1(net934),
    .B2(net867),
    .C1(net953),
    .Y(net118));
 sky130_fd_sc_hd__and2b_2 c193 (.A_N(net97),
    .B(net111),
    .X(net119));
 sky130_fd_sc_hd__a221o_2 c194 (.A1(net108),
    .A2(net118),
    .B1(net114),
    .B2(net112),
    .C1(net953),
    .X(net120));
 sky130_fd_sc_hd__a221o_1 c195 (.A1(net107),
    .A2(net117),
    .B1(net120),
    .B2(net119),
    .C1(net953),
    .X(net121));
 sky130_fd_sc_hd__a211oi_1 c196 (.A1(net102),
    .A2(net904),
    .B1(net121),
    .C1(net954),
    .Y(net122));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net114),
    .A1(net120),
    .A2(net117),
    .A3(net954),
    .S0(net121),
    .X(net123));
 sky130_fd_sc_hd__a211oi_1 c198 (.A1(net115),
    .A2(net956),
    .B1(net855),
    .C1(net867),
    .Y(net124));
 sky130_fd_sc_hd__nand3b_1 c199 (.A_N(net116),
    .B(net69),
    .C(net954),
    .Y(net125));
 sky130_fd_sc_hd__mux4_2 c200 (.A0(net847),
    .A1(net946),
    .A2(net9),
    .A3(net958),
    .S0(net125),
    .S1(net956),
    .X(net126));
 sky130_fd_sc_hd__and2_1 c201 (.A(net124),
    .B(net845),
    .X(net127));
 sky130_fd_sc_hd__and3b_1 c202 (.A_N(net862),
    .B(net12),
    .C(net956),
    .X(net128));
 sky130_fd_sc_hd__a221oi_4 c203 (.A1(net289),
    .A2(net115),
    .B1(net956),
    .B2(net21),
    .C1(net845),
    .Y(net129));
 sky130_fd_sc_hd__or3_4 c204 (.A(net125),
    .B(net0),
    .C(net830),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net128),
    .A1(net121),
    .A2(net916),
    .A3(net127),
    .S0(net126),
    .S1(net951),
    .X(net131));
 sky130_fd_sc_hd__nand2b_4 c206 (.A_N(net127),
    .B(net129),
    .Y(net132));
 sky130_fd_sc_hd__or3_2 c207 (.A(net75),
    .B(net9),
    .C(net955),
    .X(net133));
 sky130_fd_sc_hd__nand3_2 c208 (.A(net133),
    .B(net956),
    .C(net825),
    .Y(net134));
 sky130_fd_sc_hd__a211oi_2 c209 (.A1(net830),
    .A2(net129),
    .B1(net207),
    .C1(net956),
    .Y(net135));
 sky130_fd_sc_hd__or3b_4 c210 (.A(net855),
    .B(net134),
    .C_N(net956),
    .X(net876));
 sky130_fd_sc_hd__nor3_1 c211 (.A(net21),
    .B(net958),
    .C(net951),
    .Y(net136));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net121),
    .A1(net19),
    .A2(net135),
    .A3(net876),
    .S0(net956),
    .X(net137));
 sky130_fd_sc_hd__mux4_2 c213 (.A0(net134),
    .A1(net6),
    .A2(net956),
    .A3(net126),
    .S0(net876),
    .S1(net696),
    .X(net905));
 sky130_fd_sc_hd__a211o_1 c214 (.A1(net109),
    .A2(net945),
    .B1(net135),
    .C1(net696),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net135),
    .A1(net876),
    .A2(net127),
    .A3(net132),
    .S0(net133),
    .S1(net931),
    .X(net139));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net135),
    .A1(net130),
    .A2(net931),
    .A3(net957),
    .S0(net23),
    .S1(net700),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net140),
    .A1(net133),
    .A2(net126),
    .A3(net135),
    .S0(net905),
    .S1(net130),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net23),
    .A1(net133),
    .A2(net135),
    .A3(net132),
    .S0(net696),
    .S1(net735),
    .X(net142));
 sky130_fd_sc_hd__mux4_2 c219 (.A0(net136),
    .A1(net139),
    .A2(net6),
    .A3(net931),
    .S0(net134),
    .S1(net736),
    .X(net143));
 sky130_fd_sc_hd__and2b_2 c220 (.A_N(net33),
    .B(net876),
    .X(net144));
 sky130_fd_sc_hd__and3_2 c221 (.A(net19),
    .B(net36),
    .C(net28),
    .X(net922));
 sky130_fd_sc_hd__nor2b_1 c222 (.A(net118),
    .B_N(net34),
    .Y(net145));
 sky130_fd_sc_hd__nor2b_1 c223 (.A(net908),
    .B_N(net700),
    .Y(net146));
 sky130_fd_sc_hd__or3_1 c224 (.A(net69),
    .B(net822),
    .C(net931),
    .X(net147));
 sky130_fd_sc_hd__nor2_2 c225 (.A(net101),
    .B(net34),
    .Y(net892));
 sky130_fd_sc_hd__buf_2 c226 (.A(net728),
    .X(net148));
 sky130_fd_sc_hd__or2_2 c227 (.A(net29),
    .B(net736),
    .X(net149));
 sky130_fd_sc_hd__inv_4 c228 (.A(net728),
    .Y(net150));
 sky130_fd_sc_hd__inv_1 c229 (.A(net708),
    .Y(net151));
 sky130_fd_sc_hd__mux4_4 c230 (.A0(net147),
    .A1(net149),
    .A2(net25),
    .A3(net24),
    .S0(net148),
    .S1(net700),
    .X(net152));
 sky130_fd_sc_hd__a221oi_2 c231 (.A1(net861),
    .A2(net33),
    .B1(net905),
    .B2(net150),
    .C1(net931),
    .Y(net153));
 sky130_fd_sc_hd__a211oi_4 c232 (.A1(net146),
    .A2(net951),
    .B1(net931),
    .C1(net101),
    .Y(net154));
 sky130_fd_sc_hd__a221oi_1 c233 (.A1(net892),
    .A2(net931),
    .B1(net834),
    .B2(net700),
    .C1(net993),
    .Y(net155));
 sky130_fd_sc_hd__clkbuf_1 c234 (.A(net655),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 c235 (.A(net727),
    .X(net157));
 sky130_fd_sc_hd__and3b_1 c236 (.A_N(net156),
    .B(net28),
    .C(net118),
    .X(net158));
 sky130_fd_sc_hd__a221oi_1 c237 (.A1(net157),
    .A2(net158),
    .B1(net156),
    .B2(net153),
    .C1(net978),
    .Y(net159));
 sky130_fd_sc_hd__sdfbbn_2 c238 (.CLK_N(clknet_4_15_0_clk),
    .D(net157),
    .RESET_B(net138),
    .SCD(net154),
    .SCE(net158),
    .SET_B(net148),
    .Q(net161),
    .Q_N(net160));
 sky130_fd_sc_hd__a211oi_1 c239 (.A1(net151),
    .A2(net154),
    .B1(net158),
    .C1(net876),
    .Y(net162));
 sky130_fd_sc_hd__a211oi_1 c240 (.A1(net922),
    .A2(net921),
    .B1(net721),
    .C1(net919),
    .Y(net163));
 sky130_fd_sc_hd__mux4_2 c241 (.A0(net163),
    .A1(net157),
    .A2(net69),
    .A3(net905),
    .S0(net867),
    .S1(net721),
    .X(net164));
 sky130_fd_sc_hd__a211oi_1 c242 (.A1(net148),
    .A2(net905),
    .B1(net922),
    .C1(net898),
    .Y(net900));
 sky130_fd_sc_hd__a211oi_4 c243 (.A1(net35),
    .A2(net905),
    .B1(net207),
    .C1(net24),
    .Y(net165));
 sky130_fd_sc_hd__o21ba_1 c244 (.A1(net149),
    .A2(net35),
    .B1_N(net931),
    .X(net887));
 sky130_fd_sc_hd__a211oi_1 c245 (.A1(net18),
    .A2(net149),
    .B1(net47),
    .C1(net945),
    .Y(net166));
 sky130_fd_sc_hd__o21a_2 c246 (.A1(net54),
    .A2(net56),
    .B1(net945),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_1 c247 (.A(net804),
    .X(net167));
 sky130_fd_sc_hd__a211oi_1 c248 (.A1(net931),
    .A2(net837),
    .B1(net895),
    .C1(net165),
    .Y(net168));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net24),
    .A1(net910),
    .A2(net895),
    .A3(net887),
    .S0(net908),
    .S1(net919),
    .X(net169));
 sky130_fd_sc_hd__sdfrbp_1 c250 (.CLK(clknet_4_15_0_clk),
    .D(net167),
    .RESET_B(net895),
    .SCD(net138),
    .SCE(net896),
    .Q(net171),
    .Q_N(net170));
 sky130_fd_sc_hd__sdfrbp_1 c251 (.CLK(clknet_4_14_0_clk),
    .D(net58),
    .RESET_B(net889),
    .SCD(net895),
    .SCE(net896),
    .Q(net911),
    .Q_N(net172));
 sky130_fd_sc_hd__mux4_1 c252 (.A0(net166),
    .A1(net922),
    .A2(net18),
    .A3(net165),
    .S0(net692),
    .S1(net896),
    .X(net173));
 sky130_fd_sc_hd__a211oi_1 c253 (.A1(net817),
    .A2(net165),
    .B1(net734),
    .C1(net896),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 c254 (.A(net804),
    .Y(net891));
 sky130_fd_sc_hd__a21o_1 c255 (.A1(net867),
    .A2(net24),
    .B1(net919),
    .X(net175));
 sky130_fd_sc_hd__sdfrtn_1 c256 (.CLK_N(clknet_4_15_0_clk),
    .D(net62),
    .RESET_B(net895),
    .SCD(net165),
    .SCE(net734),
    .Q(net176));
 sky130_fd_sc_hd__mux2_1 c257 (.A0(net176),
    .A1(net61),
    .S(net913),
    .X(net914));
 sky130_fd_sc_hd__a221oi_4 c258 (.A1(net61),
    .A2(net176),
    .B1(net931),
    .B2(net170),
    .C1(net951),
    .Y(net923));
 sky130_fd_sc_hd__a211o_1 c259 (.A1(net153),
    .A2(net898),
    .B1(net165),
    .C1(net923),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net876),
    .A1(net904),
    .A2(net840),
    .A3(net923),
    .S0(net35),
    .S1(net1002),
    .X(net178));
 sky130_fd_sc_hd__a221o_1 c261 (.A1(net171),
    .A2(net24),
    .B1(net923),
    .B2(net951),
    .C1(net687),
    .X(net179));
 sky130_fd_sc_hd__mux4_4 c262 (.A0(net47),
    .A1(net923),
    .A2(net895),
    .A3(net908),
    .S0(net734),
    .S1(net896),
    .X(net180));
 sky130_fd_sc_hd__mux4_4 c263 (.A0(net175),
    .A1(net58),
    .A2(net923),
    .A3(net867),
    .S0(net910),
    .S1(net896),
    .X(net181));
 sky130_fd_sc_hd__mux2_1 c264 (.A0(net196),
    .A1(net197),
    .S(net815),
    .X(net182));
 sky130_fd_sc_hd__mux4_2 c265 (.A0(net199),
    .A1(net63),
    .A2(net200),
    .A3(net193),
    .S0(net195),
    .S1(net948),
    .X(net912));
 sky130_fd_sc_hd__and2_1 c266 (.A(net74),
    .B(net196),
    .X(net183));
 sky130_fd_sc_hd__a21oi_1 c267 (.A1(net182),
    .A2(net72),
    .B1(net195),
    .Y(net184));
 sky130_fd_sc_hd__o21bai_2 c268 (.A1(net183),
    .A2(net182),
    .B1_N(net198),
    .Y(net185));
 sky130_fd_sc_hd__mux4_2 c269 (.A0(net201),
    .A1(net68),
    .A2(net199),
    .A3(net1007),
    .S0(net195),
    .S1(net198),
    .X(net885));
 sky130_fd_sc_hd__mux2_1 c270 (.A0(net816),
    .A1(net184),
    .S(net182),
    .X(net186));
 sky130_fd_sc_hd__a21o_1 c271 (.A1(net885),
    .A2(net201),
    .B1(net185),
    .X(net187));
 sky130_fd_sc_hd__mux2_1 c272 (.A0(net198),
    .A1(net187),
    .S(net77),
    .X(net188));
 sky130_fd_sc_hd__o21ba_1 c273 (.A1(net197),
    .A2(net183),
    .B1_N(net82),
    .X(net189));
 sky130_fd_sc_hd__o21ba_2 c274 (.A1(net187),
    .A2(net188),
    .B1_N(net936),
    .X(net190));
 sky130_fd_sc_hd__a221o_1 c275 (.A1(net186),
    .A2(net969),
    .B1(net190),
    .B2(net936),
    .C1(net948),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c276 (.A0(net190),
    .A1(net186),
    .A2(net82),
    .A3(net187),
    .S0(net969),
    .S1(net1000),
    .X(net192));
 sky130_fd_sc_hd__and2_1 c277 (.A(net843),
    .B(net78),
    .X(net193));
 sky130_fd_sc_hd__or2_1 c278 (.A(net820),
    .B(net45),
    .X(net194));
 sky130_fd_sc_hd__and2b_2 c279 (.A_N(net78),
    .B(net72),
    .X(net195));
 sky130_fd_sc_hd__nand2_4 c280 (.A(net195),
    .B(net975),
    .Y(net196));
 sky130_fd_sc_hd__o21ai_4 c281 (.A1(net193),
    .A2(net939),
    .B1(net45),
    .Y(net197));
 sky130_fd_sc_hd__and2_1 c282 (.A(net195),
    .B(net82),
    .X(net198));
 sky130_fd_sc_hd__a21bo_2 c283 (.A1(net77),
    .A2(net198),
    .B1_N(net949),
    .X(net199));
 sky130_fd_sc_hd__a21bo_1 c284 (.A1(net197),
    .A2(net195),
    .B1_N(net947),
    .X(net200));
 sky130_fd_sc_hd__nand2_1 c285 (.A(net1007),
    .B(net872),
    .Y(net201));
 sky130_fd_sc_hd__or2_1 c286 (.A(net96),
    .B(net83),
    .X(net202));
 sky130_fd_sc_hd__or2_1 c287 (.A(net188),
    .B(net100),
    .X(net203));
 sky130_fd_sc_hd__nor2b_4 c288 (.A(net935),
    .B_N(net830),
    .Y(net204));
 sky130_fd_sc_hd__a21o_1 c289 (.A1(net83),
    .A2(net94),
    .B1(net85),
    .X(net205));
 sky130_fd_sc_hd__or2b_1 c290 (.A(net205),
    .B_N(net90),
    .X(net206));
 sky130_fd_sc_hd__inv_1 c293_4 (.A(clknet_1_1__leaf_net706),
    .Y(net962));
 sky130_fd_sc_hd__inv_4 c292 (.A(net713),
    .Y(net208));
 sky130_fd_sc_hd__inv_6 c425_8 (.A(clknet_1_1__leaf_net707),
    .Y(net966));
 sky130_fd_sc_hd__o21ai_0 c294 (.A1(net965),
    .A2(net199),
    .B1(net202),
    .Y(net210));
 sky130_fd_sc_hd__nor2_1 c295 (.A(net86),
    .B(net208),
    .Y(net211));
 sky130_fd_sc_hd__o21bai_1 c296 (.A1(net210),
    .A2(net835),
    .B1_N(net830),
    .Y(net212));
 sky130_fd_sc_hd__mux4_1 c297 (.A0(net100),
    .A1(net211),
    .A2(net206),
    .A3(net208),
    .S0(net205),
    .S1(net949),
    .X(net213));
 sky130_fd_sc_hd__a21o_2 c298 (.A1(net208),
    .A2(net188),
    .B1(net196),
    .X(net214));
 sky130_fd_sc_hd__a21o_1 c299 (.A1(net830),
    .A2(net92),
    .B1(net936),
    .X(net215));
 sky130_fd_sc_hd__a21boi_2 c300 (.A1(net825),
    .A2(net961),
    .B1_N(net205),
    .Y(net216));
 sky130_fd_sc_hd__mux4_2 c301 (.A0(net960),
    .A1(net964),
    .A2(net208),
    .A3(net204),
    .S0(net844),
    .S1(net199),
    .X(net217));
 sky130_fd_sc_hd__mux4_2 c302 (.A0(net216),
    .A1(net949),
    .A2(net215),
    .A3(net90),
    .S0(net95),
    .S1(net830),
    .X(net218));
 sky130_fd_sc_hd__mux2_4 c303 (.A0(net215),
    .A1(net963),
    .S(clknet_1_1__leaf_net218),
    .X(net219));
 sky130_fd_sc_hd__and2_1 c304 (.A(net211),
    .B(net206),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net213),
    .A1(net204),
    .A2(net208),
    .A3(net959),
    .S0(clknet_1_1__leaf_net218),
    .S1(clknet_1_1__leaf_net219),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net220),
    .A1(net83),
    .A2(net205),
    .A3(net90),
    .S0(net92),
    .S1(clknet_1_0__leaf_net706),
    .X(net222));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net222),
    .A1(net815),
    .A2(net220),
    .A3(net215),
    .S0(net832),
    .S1(clknet_1_1__leaf_net218),
    .X(net223));
 sky130_fd_sc_hd__inv_2 c308 (.A(net691),
    .Y(net224));
 sky130_fd_sc_hd__a211o_1 c309 (.A1(net848),
    .A2(net224),
    .B1(net45),
    .C1(net955),
    .X(net225));
 sky130_fd_sc_hd__o21bai_1 c310 (.A1(net941),
    .A2(net936),
    .B1_N(clknet_1_1__leaf_net706),
    .Y(net226));
 sky130_fd_sc_hd__and2b_2 c311 (.A_N(net934),
    .B(clknet_1_1__leaf_net706),
    .X(net227));
 sky130_fd_sc_hd__nor2_1 c312 (.A(net853),
    .B(net936),
    .Y(net228));
 sky130_fd_sc_hd__a21oi_4 c313 (.A1(net860),
    .A2(net841),
    .B1(net119),
    .Y(net229));
 sky130_fd_sc_hd__o21ai_1 c314 (.A1(net852),
    .A2(net106),
    .B1(net939),
    .Y(net230));
 sky130_fd_sc_hd__a21o_1 c315 (.A1(net858),
    .A2(net119),
    .B1(net958),
    .X(net231));
 sky130_fd_sc_hd__o21a_1 c316 (.A1(net228),
    .A2(net936),
    .B1(clknet_1_0__leaf_net706),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 c317 (.A(net691),
    .X(net233));
 sky130_fd_sc_hd__a21oi_2 c318 (.A1(net230),
    .A2(net233),
    .B1(clknet_1_1__leaf_net706),
    .Y(net234));
 sky130_fd_sc_hd__a21o_4 c319 (.A1(net224),
    .A2(net228),
    .B1(net955),
    .X(net893));
 sky130_fd_sc_hd__mux2_2 c320 (.A0(net941),
    .A1(net830),
    .S(net955),
    .X(net235));
 sky130_fd_sc_hd__a21bo_2 c321 (.A1(net119),
    .A2(net933),
    .B1_N(clknet_1_0__leaf_net234),
    .X(net236));
 sky130_fd_sc_hd__mux2_1 c322 (.A0(net231),
    .A1(net228),
    .S(net230),
    .X(net237));
 sky130_fd_sc_hd__a21oi_4 c323 (.A1(net226),
    .A2(net934),
    .B1(net940),
    .Y(net238));
 sky130_fd_sc_hd__nor2_2 c324 (.A(net227),
    .B(net940),
    .Y(net239));
 sky130_fd_sc_hd__a211oi_2 c325 (.A1(net233),
    .A2(net893),
    .B1(net82),
    .C1(clknet_1_0__leaf_net217),
    .Y(net240));
 sky130_fd_sc_hd__a221oi_4 c326 (.A1(net88),
    .A2(net940),
    .B1(clknet_1_1__leaf_net240),
    .B2(net835),
    .C1(net955),
    .Y(net241));
 sky130_fd_sc_hd__buf_1 c327 (.A(net713),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 c328 (.A(net807),
    .X(net899));
 sky130_fd_sc_hd__mux4_4 c329 (.A0(net938),
    .A1(clknet_1_0__leaf_net234),
    .A2(clknet_1_0__leaf_net241),
    .A3(net958),
    .S0(net940),
    .S1(clknet_1_1__leaf_net706),
    .X(net243));
 sky130_fd_sc_hd__a211oi_1 c330 (.A1(net92),
    .A2(net132),
    .B1(net242),
    .C1(net972),
    .Y(net244));
 sky130_fd_sc_hd__a21o_1 c331 (.A1(net233),
    .A2(net126),
    .B1(net204),
    .X(net245));
 sky130_fd_sc_hd__mux4_4 c332 (.A0(clknet_1_1__leaf_net217),
    .A1(net132),
    .A2(net973),
    .A3(net0),
    .S0(net957),
    .S1(net929),
    .X(net246));
 sky130_fd_sc_hd__mux2_4 c333 (.A0(net212),
    .A1(clknet_1_0__leaf_net239),
    .S(net935),
    .X(net247));
 sky130_fd_sc_hd__o21ba_1 c334 (.A1(net245),
    .A2(net126),
    .B1_N(net825),
    .X(net248));
 sky130_fd_sc_hd__a211o_1 c335 (.A1(net142),
    .A2(net12),
    .B1(net929),
    .C1(clknet_1_1__leaf_net247),
    .X(net249));
 sky130_fd_sc_hd__a21o_1 c336 (.A1(net957),
    .A2(net9),
    .B1(net940),
    .X(net250));
 sky130_fd_sc_hd__clkinv_4 c337 (.A(net805),
    .Y(net897));
 sky130_fd_sc_hd__sdfrtp_1 c338 (.CLK(clknet_4_7_0_clk),
    .D(net841),
    .RESET_B(clknet_1_1__leaf_net239),
    .SCD(net248),
    .SCE(net830),
    .Q(net251));
 sky130_fd_sc_hd__a211o_4 c339 (.A1(net251),
    .A2(net897),
    .B1(net899),
    .C1(net957),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(clknet_1_1__leaf_net247),
    .A1(net242),
    .A2(net252),
    .A3(net905),
    .S0(net929),
    .X(net253));
 sky130_fd_sc_hd__a21boi_0 c341 (.A1(clknet_1_0__leaf_net239),
    .A2(net245),
    .B1_N(net250),
    .Y(net254));
 sky130_fd_sc_hd__a221o_1 c342 (.A1(net238),
    .A2(net973),
    .B1(clknet_1_1__leaf_net254),
    .B2(net907),
    .C1(net929),
    .X(net255));
 sky130_fd_sc_hd__a21o_1 c343 (.A1(net962),
    .A2(net897),
    .B1(net132),
    .X(net256));
 sky130_fd_sc_hd__inv_4 c344 (.A(net805),
    .Y(net257));
 sky130_fd_sc_hd__sdfbbn_2 c345 (.CLK_N(clknet_4_13_0_clk),
    .D(net242),
    .RESET_B(net984),
    .SCD(net90),
    .SCE(net929),
    .SET_B(clknet_1_0__leaf_net247),
    .Q(net259),
    .Q_N(net258));
 sky130_fd_sc_hd__sdfbbp_1 c346 (.CLK(clknet_4_13_0_clk),
    .D(net126),
    .RESET_B(net929),
    .SCD(clknet_1_0__leaf_net256),
    .SCE(net258),
    .SET_B(net984),
    .Q(net261),
    .Q_N(net260));
 sky130_fd_sc_hd__a221o_1 c347 (.A1(net257),
    .A2(net258),
    .B1(net929),
    .B2(net698),
    .C1(net713),
    .X(net262));
 sky130_fd_sc_hd__a211oi_1 c348 (.A1(net261),
    .A2(net951),
    .B1(net698),
    .C1(net717),
    .Y(net263));
 sky130_fd_sc_hd__inv_4 c349 (.A(net709),
    .Y(net264));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(clknet_1_0__leaf_net247),
    .A1(net251),
    .A2(net264),
    .A3(net252),
    .S0(net258),
    .S1(net132),
    .X(net265));
 sky130_fd_sc_hd__o21ba_1 c351 (.A1(net817),
    .A2(net713),
    .B1_N(clknet_1_1__leaf_net738),
    .X(net266));
 sky130_fd_sc_hd__or2b_2 c352 (.A(net34),
    .B_N(net904),
    .X(net267));
 sky130_fd_sc_hd__nor2b_2 c353 (.A(net12),
    .B_N(net148),
    .Y(net268));
 sky130_fd_sc_hd__clkbuf_2 c354 (.A(net636),
    .X(net269));
 sky130_fd_sc_hd__and2_1 c355 (.A(net29),
    .B(net252),
    .X(net270));
 sky130_fd_sc_hd__nand2_1 c356 (.A(net268),
    .B(net908),
    .Y(net918));
 sky130_fd_sc_hd__nand2_1 c357 (.A(net270),
    .B(net899),
    .Y(net271));
 sky130_fd_sc_hd__mux4_2 c358 (.A0(net269),
    .A1(net164),
    .A2(net268),
    .A3(net937),
    .S0(net267),
    .S1(clknet_1_0__leaf_net881),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 c359 (.A(net636),
    .X(net273));
 sky130_fd_sc_hd__inv_2 c360 (.A(net656),
    .Y(net274));
 sky130_fd_sc_hd__nor2_2 c361 (.A(net273),
    .B(net269),
    .Y(net902));
 sky130_fd_sc_hd__or2_1 c362 (.A(net6),
    .B(net269),
    .X(net275));
 sky130_fd_sc_hd__nor2b_1 c363 (.A(net271),
    .B_N(net976),
    .Y(net276));
 sky130_fd_sc_hd__mux4_4 c364 (.A0(net267),
    .A1(net275),
    .A2(net269),
    .A3(net271),
    .S0(net148),
    .S1(clknet_1_0__leaf_net881),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net274),
    .A1(net267),
    .A2(net276),
    .A3(net922),
    .S0(net12),
    .S1(net940),
    .X(net278));
 sky130_fd_sc_hd__mux4_4 c366 (.A0(net275),
    .A1(net161),
    .A2(net267),
    .A3(net897),
    .S0(net269),
    .S1(clknet_1_1__leaf_net739),
    .X(net279));
 sky130_fd_sc_hd__or2_1 c367 (.A(net908),
    .B(net697),
    .X(net280));
 sky130_fd_sc_hd__mux4_4 c368 (.A0(net2),
    .A1(net269),
    .A2(clknet_1_1__leaf_net256),
    .A3(clknet_1_1__leaf_net739),
    .S0(net740),
    .S1(net743),
    .X(net281));
 sky130_fd_sc_hd__nand2_1 c369 (.A(net276),
    .B(net252),
    .Y(net282));
 sky130_fd_sc_hd__mux4_4 c370 (.A0(net9),
    .A1(clknet_1_1__leaf_net256),
    .A2(net12),
    .A3(net740),
    .S0(net742),
    .S1(net744),
    .X(net283));
 sky130_fd_sc_hd__and2_2 c371 (.A(net37),
    .B(net275),
    .X(net284));
 sky130_fd_sc_hd__mux4_2 c372 (.A0(net284),
    .A1(net280),
    .A2(net894),
    .A3(clknet_1_1__leaf_net881),
    .S0(net743),
    .S1(net744),
    .X(net285));
 sky130_fd_sc_hd__mux4_2 c373 (.A0(net158),
    .A1(net280),
    .A2(net973),
    .A3(net284),
    .S0(net268),
    .S1(net742),
    .X(net286));
 sky130_fd_sc_hd__mux4_2 c392 (.A0(net282),
    .A1(net897),
    .A2(net172),
    .A3(net908),
    .S0(net917),
    .S1(net896),
    .X(net920));
 sky130_fd_sc_hd__mux4_4 c393 (.A0(net280),
    .A1(net979),
    .A2(net920),
    .A3(net45),
    .S0(net282),
    .S1(net908),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net920),
    .A1(net282),
    .A2(net1006),
    .A3(net721),
    .S0(net990),
    .S1(net915),
    .X(net288));
 sky130_fd_sc_hd__mux4_2 c395 (.A0(net285),
    .A1(net910),
    .A2(net920),
    .A3(net892),
    .S1(net915),
    .X(net879));
 sky130_fd_sc_hd__nor2_2 c396 (.A(net75),
    .B(net81),
    .Y(net290));
 sky130_fd_sc_hd__nor2_2 c397 (.A(net185),
    .B(net1000),
    .Y(net291));
 sky130_fd_sc_hd__nor2_1 c398 (.A(net185),
    .B(net290),
    .Y(net292));
 sky130_fd_sc_hd__and2_1 c399 (.A(net290),
    .B(net935),
    .X(net293));
 sky130_fd_sc_hd__a21boi_2 c400 (.A1(net63),
    .A2(net291),
    .B1_N(net81),
    .Y(net294));
 sky130_fd_sc_hd__nor2_4 c401 (.A(net813),
    .B(net868),
    .Y(net295));
 sky130_fd_sc_hd__mux4_2 c402 (.A0(net868),
    .A1(net939),
    .A2(net63),
    .A3(net294),
    .S0(net290),
    .S1(net295),
    .X(net296));
 sky130_fd_sc_hd__nand2_4 c403 (.A(net70),
    .B(net947),
    .Y(net297));
 sky130_fd_sc_hd__nor2_4 c404 (.A(net296),
    .B(net294),
    .Y(net298));
 sky130_fd_sc_hd__o21ba_1 c405 (.A1(net865),
    .A2(net868),
    .B1_N(net295),
    .X(net299));
 sky130_fd_sc_hd__o21a_2 c406 (.A1(net292),
    .A2(net296),
    .B1(net290),
    .X(net300));
 sky130_fd_sc_hd__a221oi_1 c407 (.A1(net295),
    .A2(net294),
    .B1(net292),
    .B2(net300),
    .C1(net298),
    .Y(net301));
 sky130_fd_sc_hd__buf_4 c408 (.A(net689),
    .X(net302));
 sky130_fd_sc_hd__sdfbbn_1 c409 (.CLK_N(clknet_4_5_0_clk),
    .D(net82),
    .RESET_B(net302),
    .SCD(net290),
    .SCE(net300),
    .SET_B(net291),
    .Q(net304),
    .Q_N(net303));
 sky130_fd_sc_hd__o21bai_2 c410 (.A1(net304),
    .A2(net293),
    .B1_N(net689),
    .Y(net305));
 sky130_fd_sc_hd__o21ai_1 c411 (.A1(net302),
    .A2(net297),
    .B1(net304),
    .Y(net306));
 sky130_fd_sc_hd__a21bo_1 c412 (.A1(net305),
    .A2(net199),
    .B1_N(net292),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 c413 (.A(net689),
    .X(net308));
 sky130_fd_sc_hd__a221o_1 c414 (.A1(net306),
    .A2(net291),
    .B1(net308),
    .B2(net303),
    .C1(net947),
    .X(net309));
 sky130_fd_sc_hd__mux4_4 c415 (.A0(net294),
    .A1(net198),
    .A2(net296),
    .A3(net302),
    .S0(net300),
    .S1(net308),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net307),
    .A1(net309),
    .A2(net190),
    .A3(net950),
    .S0(net688),
    .S1(net746),
    .X(net311));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net308),
    .A1(net307),
    .A2(net305),
    .A3(net293),
    .S0(net296),
    .S1(net747),
    .X(net312));
 sky130_fd_sc_hd__inv_2 c418 (.A(net720),
    .Y(net313));
 sky130_fd_sc_hd__a21oi_1 c419 (.A1(net94),
    .A2(net843),
    .B1(net747),
    .Y(net314));
 sky130_fd_sc_hd__or2b_4 c420 (.A(net843),
    .B_N(net290),
    .X(net315));
 sky130_fd_sc_hd__o21bai_1 c421 (.A1(net208),
    .A2(net309),
    .B1_N(net299),
    .Y(net316));
 sky130_fd_sc_hd__and2_0 c422 (.A(net936),
    .B(net75),
    .X(net317));
 sky130_fd_sc_hd__buf_12 c423 (.A(clknet_1_0__leaf_net707),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 c424 (.A(net720),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__and2_2 c426 (.A(net293),
    .B(net75),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c427 (.A0(net316),
    .A1(net204),
    .A2(net844),
    .A3(net297),
    .S0(clknet_1_1__leaf_net219),
    .S1(net746),
    .X(net322));
 sky130_fd_sc_hd__a211oi_1 c428 (.A1(net203),
    .A2(net319),
    .B1(net84),
    .C1(net1003),
    .Y(net323));
 sky130_fd_sc_hd__sdfbbn_1 c429 (.CLK_N(clknet_4_5_0_clk),
    .D(net321),
    .RESET_B(net315),
    .SCD(net214),
    .SCE(net293),
    .SET_B(net670),
    .Q(net325),
    .Q_N(net324));
 sky130_fd_sc_hd__sdfrtp_4 c430 (.CLK(clknet_4_5_0_clk),
    .D(net844),
    .RESET_B(net214),
    .SCD(net314),
    .SCE(net670),
    .Q(net326));
 sky130_fd_sc_hd__or2_1 c431 (.A(net309),
    .B(net835),
    .X(net327));
 sky130_fd_sc_hd__a221oi_1 c432 (.A1(net313),
    .A2(net315),
    .B1(net326),
    .B2(net297),
    .C1(net316),
    .Y(net328));
 sky130_fd_sc_hd__a211oi_4 c433 (.A1(net326),
    .A2(clknet_1_0__leaf_net217),
    .B1(net321),
    .C1(net747),
    .Y(net329));
 sky130_fd_sc_hd__a21o_4 c434 (.A1(net299),
    .A2(clknet_1_0__leaf_net329),
    .B1(net746),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net318),
    .A1(net68),
    .A2(clknet_1_0__leaf_net218),
    .A3(net290),
    .S0(net315),
    .S1(net746),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net319),
    .A1(net325),
    .A2(clknet_1_0__leaf_net329),
    .A3(net326),
    .S0(clknet_1_0__leaf_net331),
    .S1(net746),
    .X(net332));
 sky130_fd_sc_hd__mux4_4 c437 (.A0(net87),
    .A1(net299),
    .A2(clknet_1_0__leaf_net330),
    .A3(net821),
    .S0(net746),
    .S1(net748),
    .X(net333));
 sky130_fd_sc_hd__mux4_2 c438 (.A0(net206),
    .A1(clknet_1_0__leaf_net331),
    .A2(net325),
    .A3(net321),
    .S0(clknet_1_0__leaf_net707),
    .S1(net748),
    .X(net334));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net326),
    .A1(clknet_1_0__leaf_net331),
    .A2(net298),
    .A3(clknet_1_0__leaf_net707),
    .S0(net748),
    .S1(net749),
    .X(net335));
 sky130_fd_sc_hd__nand2b_1 c440 (.A_N(net958),
    .B(net225),
    .Y(net336));
 sky130_fd_sc_hd__sdfrtp_4 c441 (.CLK(clknet_4_7_0_clk),
    .D(net312),
    .RESET_B(net967),
    .SCD(net815),
    .SCE(net690),
    .Q(net337));
 sky130_fd_sc_hd__a21bo_1 c442 (.A1(net947),
    .A2(net327),
    .B1_N(net749),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net337),
    .A1(net832),
    .A2(net936),
    .A3(net326),
    .S0(net120),
    .S1(net312),
    .X(net339));
 sky130_fd_sc_hd__a21o_1 c444 (.A1(net326),
    .A2(net225),
    .B1(net337),
    .X(net340));
 sky130_fd_sc_hd__a21o_2 c445 (.A1(clknet_1_0__leaf_net240),
    .A2(net336),
    .B1(net947),
    .X(net341));
 sky130_fd_sc_hd__and2b_2 c446 (.A_N(net325),
    .B(clknet_1_0__leaf_net240),
    .X(net342));
 sky130_fd_sc_hd__buf_1 c447 (.A(net712),
    .X(net343));
 sky130_fd_sc_hd__a21boi_1 c448 (.A1(net327),
    .A2(net343),
    .B1_N(clknet_1_0__leaf_net329),
    .Y(net344));
 sky130_fd_sc_hd__a221o_2 c449 (.A1(net120),
    .A2(net343),
    .B1(net315),
    .B2(clknet_1_0__leaf_net342),
    .C1(clknet_1_0__leaf_net330),
    .X(net345));
 sky130_fd_sc_hd__sdfsbp_1 c450 (.CLK(clknet_4_7_0_clk),
    .D(net224),
    .SCD(net337),
    .SCE(net315),
    .SET_B(clknet_1_0__leaf_net344),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__o21bai_1 c451 (.A1(net120),
    .A2(net936),
    .B1_N(net681),
    .Y(net348));
 sky130_fd_sc_hd__mux2_1 c452 (.A0(net343),
    .A1(net690),
    .S(net719),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 c453 (.A(net712),
    .X(net350));
 sky130_fd_sc_hd__sdfbbp_1 c454 (.CLK(clknet_4_7_0_clk),
    .D(net350),
    .RESET_B(net312),
    .SCD(net337),
    .SCE(net194),
    .SET_B(clknet_1_0__leaf_net330),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__mux4_2 c455 (.A0(net348),
    .A1(net336),
    .A2(clknet_1_0__leaf_net344),
    .A3(net45),
    .S0(net690),
    .S1(net719),
    .X(net353));
 sky130_fd_sc_hd__sdfsbp_1 c456 (.CLK(clknet_4_6_0_clk),
    .D(net317),
    .SCD(net352),
    .SCE(net943),
    .SET_B(net883),
    .Q(net355),
    .Q_N(net354));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net337),
    .A1(net324),
    .A2(net936),
    .A3(net312),
    .S0(net1001),
    .S1(net349),
    .X(net356));
 sky130_fd_sc_hd__mux4_2 c458 (.A0(clknet_1_1__leaf_net331),
    .A1(net352),
    .A2(net355),
    .A3(net315),
    .S0(net302),
    .S1(net754),
    .X(net357));
 sky130_fd_sc_hd__mux2_4 c459 (.A0(net225),
    .A1(clknet_1_1__leaf_net329),
    .S(net754),
    .X(net358));
 sky130_fd_sc_hd__a211o_4 c460 (.A1(clknet_1_1__leaf_net232),
    .A2(clknet_1_1__leaf_net331),
    .B1(net893),
    .C1(net754),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net204),
    .A1(clknet_1_1__leaf_net358),
    .A2(net893),
    .A3(net883),
    .S0(net337),
    .S1(net349),
    .X(net360));
 sky130_fd_sc_hd__o21ai_1 c462 (.A1(net263),
    .A2(net302),
    .B1(net130),
    .Y(net361));
 sky130_fd_sc_hd__inv_2 c463 (.A(net644),
    .Y(net362));
 sky130_fd_sc_hd__inv_4 c464 (.A(net643),
    .Y(net363));
 sky130_fd_sc_hd__a221oi_4 c465 (.A1(net250),
    .A2(net929),
    .B1(clknet_1_1__leaf_net344),
    .B2(net977),
    .C1(net696),
    .Y(net364));
 sky130_fd_sc_hd__sdfbbn_2 c466 (.CLK_N(clknet_4_9_0_clk),
    .D(net929),
    .RESET_B(net263),
    .SCD(net945),
    .SCE(net264),
    .SET_B(net958),
    .Q(net366),
    .Q_N(net365));
 sky130_fd_sc_hd__a221o_4 c467 (.A1(net257),
    .A2(net363),
    .B1(net4),
    .B2(clknet_1_0__leaf_net881),
    .C1(net755),
    .X(net367));
 sky130_fd_sc_hd__a211o_4 c468 (.A1(clknet_1_1__leaf_net217),
    .A2(net832),
    .B1(net696),
    .C1(net755),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(clknet_1_1__leaf_net266),
    .A1(net973),
    .A2(net264),
    .A3(net132),
    .S0(net365),
    .S1(clknet_1_1__leaf_net330),
    .X(net369));
 sky130_fd_sc_hd__a211oi_2 c470 (.A1(clknet_1_1__leaf_net368),
    .A2(clknet_1_0__leaf_net266),
    .B1(net691),
    .C1(net944),
    .Y(net370));
 sky130_fd_sc_hd__a211o_1 c471 (.A1(net835),
    .A2(net363),
    .B1(net945),
    .C1(net944),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 c472 (.A(net809),
    .X(net372));
 sky130_fd_sc_hd__sdfstp_1 c473 (.CLK(clknet_4_12_0_clk),
    .D(net5),
    .SCD(clknet_1_1__leaf_net330),
    .SCE(net130),
    .SET_B(clknet_1_1__leaf_net344),
    .Q(net373));
 sky130_fd_sc_hd__sdfbbn_1 c474 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net367),
    .RESET_B(clknet_1_0__leaf_net368),
    .SCD(net366),
    .SCE(net929),
    .SET_B(net371),
    .Q(net375),
    .Q_N(net374));
 sky130_fd_sc_hd__a21oi_2 c475 (.A1(net132),
    .A2(net130),
    .B1(net371),
    .Y(net376));
 sky130_fd_sc_hd__a211o_1 c476 (.A1(net373),
    .A2(net885),
    .B1(net752),
    .C1(net755),
    .X(net377));
 sky130_fd_sc_hd__inv_2 c477 (.A(net810),
    .Y(net901));
 sky130_fd_sc_hd__sdfstp_1 c478 (.CLK(clknet_4_12_0_clk),
    .D(net372),
    .SCD(net363),
    .SCE(clknet_1_1__leaf_net330),
    .SET_B(net712),
    .Q(net378));
 sky130_fd_sc_hd__mux4_2 c479 (.A0(net362),
    .A1(clknet_1_0__leaf_net368),
    .A2(net377),
    .A3(net378),
    .S0(net374),
    .S1(clknet_1_1__leaf_net342),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net336),
    .A1(net371),
    .A2(net375),
    .A3(clknet_1_0__leaf_net368),
    .S0(net365),
    .S1(net362),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 c481 (.A(net709),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net343),
    .A1(net380),
    .A2(net5),
    .A3(net376),
    .S0(clknet_1_1__leaf_net370),
    .S1(net204),
    .X(net382));
 sky130_fd_sc_hd__mux4_4 c483 (.A0(net264),
    .A1(net381),
    .A2(clknet_1_1__leaf_net370),
    .A3(clknet_1_1__leaf_net234),
    .S0(net958),
    .S1(clknet_1_0__leaf_net757),
    .X(net383));
 sky130_fd_sc_hd__a221oi_2 c484 (.A1(net940),
    .A2(net252),
    .B1(net26),
    .B2(net680),
    .C1(net755),
    .Y(net384));
 sky130_fd_sc_hd__a221oi_4 c485 (.A1(net144),
    .A2(net366),
    .B1(net905),
    .B2(net958),
    .C1(net897),
    .Y(net385));
 sky130_fd_sc_hd__sdfbbp_1 c486 (.CLK(clknet_4_14_0_clk),
    .D(net268),
    .RESET_B(net25),
    .SCD(net385),
    .SCE(clknet_1_1__leaf_net330),
    .SET_B(net741),
    .Q(net387),
    .Q_N(net386));
 sky130_fd_sc_hd__sdfstp_1 c487 (.CLK(clknet_4_12_0_clk),
    .D(net36),
    .SCD(net975),
    .SCE(net286),
    .SET_B(net741),
    .Q(net388));
 sky130_fd_sc_hd__a221oi_2 c488 (.A1(net0),
    .A2(net902),
    .B1(net899),
    .B2(net979),
    .C1(net883),
    .Y(net389));
 sky130_fd_sc_hd__a211oi_1 c489 (.A1(net387),
    .A2(net384),
    .B1(net958),
    .C1(net985),
    .Y(net390));
 sky130_fd_sc_hd__a221o_4 c490 (.A1(net259),
    .A2(net388),
    .B1(net901),
    .B2(net375),
    .C1(net755),
    .X(net874));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net375),
    .A1(net25),
    .A2(net385),
    .A3(net384),
    .S0(net940),
    .S1(net995),
    .X(net391));
 sky130_fd_sc_hd__a221o_1 c492 (.A1(net384),
    .A2(net252),
    .B1(net897),
    .B2(net386),
    .C1(net683),
    .X(net392));
 sky130_fd_sc_hd__a221oi_1 c493 (.A1(net385),
    .A2(net874),
    .B1(net366),
    .B2(net737),
    .C1(net741),
    .Y(net393));
 sky130_fd_sc_hd__a221oi_4 c494 (.A1(clknet_1_0__leaf_net368),
    .A2(net390),
    .B1(net144),
    .B2(net374),
    .C1(clknet_1_0__leaf_net234),
    .Y(net394));
 sky130_fd_sc_hd__mux4_2 c495 (.A0(clknet_1_1__leaf_net330),
    .A1(net148),
    .A2(net259),
    .A3(clknet_1_1__leaf_net394),
    .S0(net980),
    .S1(net832),
    .X(net395));
 sky130_fd_sc_hd__a221o_1 c496 (.A1(net235),
    .A2(net259),
    .B1(net144),
    .B2(net899),
    .C1(clknet_1_0__leaf_net886),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net902),
    .A1(net385),
    .A2(net874),
    .A3(clknet_1_1__leaf_net881),
    .S0(net745),
    .S1(net755),
    .X(net397));
 sky130_fd_sc_hd__a221oi_4 c498 (.A1(net315),
    .A2(net366),
    .B1(net927),
    .B2(net144),
    .C1(net388),
    .Y(net398));
 sky130_fd_sc_hd__a221o_4 c499 (.A1(net268),
    .A2(net392),
    .B1(net398),
    .B2(clknet_1_1__leaf_net396),
    .C1(net740),
    .X(net399));
 sky130_fd_sc_hd__mux4_2 c500 (.A0(net25),
    .A1(net398),
    .A2(clknet_1_0__leaf_net399),
    .A3(net385),
    .S0(clknet_1_1__leaf_net396),
    .S1(net26),
    .X(net400));
 sky130_fd_sc_hd__a221o_2 c501 (.A1(net398),
    .A2(net259),
    .B1(clknet_1_1__leaf_net396),
    .B2(net944),
    .C1(clknet_1_0__leaf_net886),
    .X(net401));
 sky130_fd_sc_hd__a211oi_1 c502 (.A1(net398),
    .A2(net897),
    .B1(net890),
    .C1(net737),
    .Y(net875));
 sky130_fd_sc_hd__a221o_4 c503 (.A1(net958),
    .A2(net144),
    .B1(net734),
    .B2(net744),
    .C1(clknet_1_1__leaf_net886),
    .X(net402));
 sky130_fd_sc_hd__mux4_2 c504 (.A0(clknet_1_1__leaf_net399),
    .A1(net402),
    .A2(net398),
    .A3(net258),
    .S0(net927),
    .S1(net745),
    .X(net403));
 sky130_fd_sc_hd__mux4_4 c505 (.A0(net403),
    .A1(net25),
    .A2(clknet_1_0__leaf_net399),
    .A3(net26),
    .S0(net745),
    .S1(net944),
    .X(net404));
 sky130_fd_sc_hd__buf_1 c528 (.A(net722),
    .X(net405));
 sky130_fd_sc_hd__and2b_2 c529 (.A_N(net81),
    .B(net291),
    .X(net406));
 sky130_fd_sc_hd__nor2b_2 c530 (.A(net81),
    .B_N(net297),
    .Y(net407));
 sky130_fd_sc_hd__clkinv_4 c531 (.A(net694),
    .Y(net408));
 sky130_fd_sc_hd__nor2b_2 c532 (.A(net406),
    .B_N(net815),
    .Y(net409));
 sky130_fd_sc_hd__a21o_2 c533 (.A1(net193),
    .A2(net408),
    .B1(net291),
    .X(net410));
 sky130_fd_sc_hd__nand2b_2 c534 (.A_N(net406),
    .B(net713),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 c535 (.A(net722),
    .Y(net412));
 sky130_fd_sc_hd__a221o_1 c536 (.A1(net412),
    .A2(net409),
    .B1(net305),
    .B2(net411),
    .C1(net295),
    .X(net413));
 sky130_fd_sc_hd__dfbbn_2 c537 (.CLK_N(clknet_4_4_0_clk),
    .D(net999),
    .RESET_B(net413),
    .SET_B(net713),
    .Q(net415),
    .Q_N(net414));
 sky130_fd_sc_hd__a221oi_4 c538 (.A1(net411),
    .A2(net415),
    .B1(net81),
    .B2(net410),
    .C1(net295),
    .Y(net416));
 sky130_fd_sc_hd__nor2_1 c539 (.A(net305),
    .B(net406),
    .Y(net417));
 sky130_fd_sc_hd__clkbuf_1 c540 (.A(net694),
    .X(net418));
 sky130_fd_sc_hd__a211o_1 c541 (.A1(net295),
    .A2(net411),
    .B1(net989),
    .C1(net747),
    .X(net419));
 sky130_fd_sc_hd__sdfbbn_2 c542 (.CLK_N(clknet_4_1_0_clk),
    .D(net419),
    .RESET_B(net409),
    .SCD(net416),
    .SCE(net300),
    .SET_B(net988),
    .Q(net873),
    .Q_N(net420));
 sky130_fd_sc_hd__nor2_1 c543 (.A(net291),
    .B(net713),
    .Y(net421));
 sky130_fd_sc_hd__or2b_2 c544 (.A(net411),
    .B_N(net688),
    .X(net422));
 sky130_fd_sc_hd__mux2_1 c545 (.A0(net418),
    .A1(net417),
    .S(net410),
    .X(net423));
 sky130_fd_sc_hd__inv_4 c546 (.A(net694),
    .Y(net424));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(net423),
    .A1(net424),
    .A2(net408),
    .A3(net295),
    .S0(net298),
    .S1(net418),
    .X(net425));
 sky130_fd_sc_hd__mux4_4 c548 (.A0(net184),
    .A1(net405),
    .A2(net422),
    .A3(net411),
    .S0(net419),
    .S1(net760),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net405),
    .A1(net422),
    .A2(net424),
    .A3(net411),
    .S0(net420),
    .S1(net761),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 c550 (.A(net710),
    .X(net428));
 sky130_fd_sc_hd__sedfxbp_2 c551 (.CLK(clknet_4_1_0_clk),
    .D(net68),
    .DE(net408),
    .SCD(net947),
    .SCE(clknet_1_0__leaf_net330),
    .Q(net430),
    .Q_N(net429));
 sky130_fd_sc_hd__a21boi_4 c552 (.A1(net196),
    .A2(net747),
    .B1_N(net749),
    .Y(net431));
 sky130_fd_sc_hd__o21a_4 c553 (.A1(net428),
    .A2(clknet_1_0__leaf_net329),
    .B1(net821),
    .X(net432));
 sky130_fd_sc_hd__buf_1 c554 (.A(net710),
    .X(net433));
 sky130_fd_sc_hd__and2b_1 c555 (.A_N(net669),
    .B(net749),
    .X(net434));
 sky130_fd_sc_hd__a211o_1 c556 (.A1(net405),
    .A2(net298),
    .B1(net434),
    .C1(net95),
    .X(net435));
 sky130_fd_sc_hd__sedfxbp_2 c557 (.CLK(clknet_4_4_0_clk),
    .D(net328),
    .DE(net428),
    .SCD(net409),
    .SCE(net763),
    .Q(net437),
    .Q_N(net436));
 sky130_fd_sc_hd__a211o_2 c558 (.A1(net297),
    .A2(net437),
    .B1(net433),
    .C1(net749),
    .X(net438));
 sky130_fd_sc_hd__a221oi_4 c559 (.A1(net321),
    .A2(net437),
    .B1(net821),
    .B2(net196),
    .C1(net950),
    .Y(net928));
 sky130_fd_sc_hd__o21ba_2 c560 (.A1(clknet_1_0__leaf_net217),
    .A2(net437),
    .B1_N(net431),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net63),
    .A1(clknet_1_1__leaf_net439),
    .A2(clknet_1_0__leaf_net217),
    .A3(net436),
    .S0(clknet_1_0__leaf_net432),
    .S1(net747),
    .X(net440));
 sky130_fd_sc_hd__mux4_2 c562 (.A0(net438),
    .A1(net406),
    .A2(net428),
    .A3(net436),
    .S0(net669),
    .S1(net760),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(net415),
    .A1(net433),
    .A2(net928),
    .A3(net424),
    .S0(net749),
    .S1(net765),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net844),
    .A1(net442),
    .A2(net438),
    .A3(net441),
    .S0(net436),
    .S1(clknet_1_0__leaf_net330),
    .X(net443));
 sky130_fd_sc_hd__inv_2 c565 (.A(net694),
    .Y(net444));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net424),
    .A1(net444),
    .A2(net442),
    .A3(net438),
    .S0(net441),
    .S1(net414),
    .X(net445));
 sky130_fd_sc_hd__a211o_1 c567 (.A1(net321),
    .A2(net434),
    .B1(net63),
    .C1(net711),
    .X(net446));
 sky130_fd_sc_hd__mux4_2 c568 (.A0(net937),
    .A1(clknet_1_0__leaf_net329),
    .A2(net436),
    .A3(net711),
    .S0(net730),
    .S1(net759),
    .X(net447));
 sky130_fd_sc_hd__a211o_1 c569 (.A1(clknet_1_0__leaf_net439),
    .A2(net422),
    .B1(clknet_1_1__leaf_net447),
    .C1(net747),
    .X(net448));
 sky130_fd_sc_hd__mux4_2 c570 (.A0(net433),
    .A1(net446),
    .A2(net437),
    .A3(net441),
    .S0(net424),
    .S1(net765),
    .X(net449));
 sky130_fd_sc_hd__mux4_4 c571 (.A0(net438),
    .A1(net437),
    .A2(clknet_1_0__leaf_net329),
    .A3(net449),
    .S0(net730),
    .S1(net765),
    .X(net450));
 sky130_fd_sc_hd__nor2_4 c572 (.A(net409),
    .B(net431),
    .Y(net451));
 sky130_fd_sc_hd__sdfbbn_1 c573 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net232),
    .RESET_B(net989),
    .SCD(net229),
    .SCE(clknet_1_0__leaf_net432),
    .SET_B(net764),
    .Q(net453),
    .Q_N(net452));
 sky130_fd_sc_hd__a211o_2 c574 (.A1(net453),
    .A2(clknet_1_0__leaf_net232),
    .B1(net893),
    .C1(net753),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 c575 (.A(net650),
    .X(net455));
 sky130_fd_sc_hd__nor2_4 c576 (.A(clknet_1_1__leaf_net454),
    .B(net766),
    .Y(net456));
 sky130_fd_sc_hd__clkbuf_1 c577 (.A(net649),
    .X(net457));
 sky130_fd_sc_hd__sedfxtp_1 c578 (.CLK(clknet_4_6_0_clk),
    .D(net355),
    .DE(net229),
    .SCD(net452),
    .SCE(clknet_1_0__leaf_net330),
    .Q(net458));
 sky130_fd_sc_hd__a21o_1 c579 (.A1(net229),
    .A2(net340),
    .B1(net766),
    .X(net459));
 sky130_fd_sc_hd__buf_1 c580 (.A(net808),
    .X(net460));
 sky130_fd_sc_hd__a221o_1 c581 (.A1(net457),
    .A2(net302),
    .B1(net460),
    .B2(net340),
    .C1(net750),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net415),
    .A1(net434),
    .A2(net461),
    .A3(net406),
    .S0(net935),
    .S1(net942),
    .X(net462));
 sky130_fd_sc_hd__mux2_4 c583 (.A0(net461),
    .A1(net457),
    .S(net459),
    .X(net463));
 sky130_fd_sc_hd__sdfbbp_1 c584 (.CLK(clknet_4_3_0_clk),
    .D(net408),
    .RESET_B(net451),
    .SCD(net459),
    .SCE(clknet_1_0__leaf_net454),
    .SET_B(net463),
    .Q(net465),
    .Q_N(net464));
 sky130_fd_sc_hd__o21ba_2 c585 (.A1(net460),
    .A2(net461),
    .B1_N(net414),
    .X(net882));
 sky130_fd_sc_hd__sdfbbn_1 c586 (.CLK_N(clknet_4_3_0_clk),
    .D(net441),
    .RESET_B(net229),
    .SCD(net882),
    .SCE(net459),
    .SET_B(net451),
    .Q(net467),
    .Q_N(net466));
 sky130_fd_sc_hd__mux4_4 c587 (.A0(net455),
    .A1(net459),
    .A2(net312),
    .A3(clknet_1_0__leaf_net454),
    .S0(clknet_1_0__leaf_net219),
    .S1(net763),
    .X(net468));
 sky130_fd_sc_hd__a21oi_1 c588 (.A1(net462),
    .A2(net453),
    .B1(net930),
    .Y(net469));
 sky130_fd_sc_hd__sdfbbn_1 c589 (.CLK_N(clknet_4_3_0_clk),
    .D(net465),
    .RESET_B(net463),
    .SCD(net882),
    .SCE(clknet_1_0__leaf_net330),
    .SET_B(net674),
    .Q(net471),
    .Q_N(net470));
 sky130_fd_sc_hd__sedfxtp_4 c590 (.CLK(clknet_4_3_0_clk),
    .D(net347),
    .DE(net469),
    .SCD(net229),
    .SCE(net409),
    .Q(net472));
 sky130_fd_sc_hd__mux4_4 c591 (.A0(net406),
    .A1(net95),
    .A2(net453),
    .A3(net459),
    .S0(net992),
    .S1(net451),
    .X(net473));
 sky130_fd_sc_hd__sdfbbp_1 c592 (.CLK(clknet_4_3_0_clk),
    .D(net467),
    .RESET_B(net459),
    .SCD(net463),
    .SCE(net312),
    .SET_B(net414),
    .Q(net878),
    .Q_N(net474));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net469),
    .A1(net470),
    .A2(clknet_1_0__leaf_net234),
    .A3(net474),
    .S0(net466),
    .S1(net674),
    .X(net475));
 sky130_fd_sc_hd__a21bo_1 c594 (.A1(net438),
    .A2(net815),
    .B1_N(net933),
    .X(net476));
 sky130_fd_sc_hd__a21boi_4 c595 (.A1(net815),
    .A2(net937),
    .B1_N(net1004),
    .Y(net477));
 sky130_fd_sc_hd__a21boi_1 c596 (.A1(net361),
    .A2(net817),
    .B1_N(net477),
    .Y(net478));
 sky130_fd_sc_hd__a221o_2 c597 (.A1(clknet_1_0__leaf_net456),
    .A2(net873),
    .B1(net324),
    .B2(net477),
    .C1(net753),
    .X(net479));
 sky130_fd_sc_hd__sdfbbn_1 c598 (.CLK_N(clknet_4_3_0_clk),
    .D(net340),
    .RESET_B(net422),
    .SCD(net431),
    .SCE(net458),
    .SET_B(net472),
    .Q(net903),
    .Q_N(net480));
 sky130_fd_sc_hd__clkbuf_2 c599 (.A(net803),
    .X(net481));
 sky130_fd_sc_hd__inv_1 c600 (.A(net803),
    .Y(net482));
 sky130_fd_sc_hd__a211o_2 c601 (.A1(net458),
    .A2(net476),
    .B1(net361),
    .C1(net716),
    .X(net884));
 sky130_fd_sc_hd__dlymetal6s2s_1 c602 (.A(net806),
    .X(net483));
 sky130_fd_sc_hd__sdfbbn_2 c603 (.CLK_N(clknet_4_6_0_clk),
    .D(net130),
    .RESET_B(clknet_1_1__leaf_net479),
    .SCD(net422),
    .SCE(net451),
    .SET_B(net716),
    .Q(net485),
    .Q_N(net484));
 sky130_fd_sc_hd__mux4_4 c604 (.A0(net422),
    .A1(net480),
    .A2(net347),
    .A3(net477),
    .S0(net481),
    .S1(net951),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_1__leaf_net342),
    .A1(net483),
    .A2(net485),
    .A3(net943),
    .S0(clknet_1_0__leaf_net370),
    .S1(clknet_1_0__leaf_net758),
    .X(net487));
 sky130_fd_sc_hd__a221oi_4 c606 (.A1(net943),
    .A2(net893),
    .B1(net933),
    .B2(clknet_1_0__leaf_net758),
    .C1(net768),
    .Y(net488));
 sky130_fd_sc_hd__mux4_2 c607 (.A0(net481),
    .A1(net438),
    .A2(clknet_1_1__leaf_net488),
    .A3(net420),
    .S0(net484),
    .S1(clknet_1_1__leaf_net758),
    .X(net489));
 sky130_fd_sc_hd__buf_1 c608 (.A(net806),
    .X(net490));
 sky130_fd_sc_hd__a21o_2 c609 (.A1(net483),
    .A2(net482),
    .B1(net481),
    .X(net491));
 sky130_fd_sc_hd__mux4_2 c610 (.A0(clknet_1_0__leaf_net488),
    .A1(net483),
    .A2(net485),
    .A3(net817),
    .S0(clknet_1_0__leaf_net489),
    .S1(net431),
    .X(net492));
 sky130_fd_sc_hd__a21boi_4 c611 (.A1(net490),
    .A2(clknet_1_1__leaf_net489),
    .B1_N(clknet_1_0__leaf_net881),
    .Y(net493));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net478),
    .A1(net491),
    .A2(clknet_1_1__leaf_net489),
    .A3(net477),
    .S1(net763),
    .X(net494));
 sky130_fd_sc_hd__a221o_1 c613 (.A1(net434),
    .A2(net252),
    .B1(net476),
    .B2(net695),
    .C1(net767),
    .X(net495));
 sky130_fd_sc_hd__mux4_4 c614 (.A0(net495),
    .A1(net491),
    .A2(net873),
    .A3(net480),
    .S0(net483),
    .S1(net87),
    .X(net496));
 sky130_fd_sc_hd__sdfbbp_1 c615 (.CLK(clknet_4_8_0_clk),
    .D(net496),
    .RESET_B(clknet_1_1__leaf_net432),
    .SCD(net490),
    .SCE(clknet_1_1__leaf_net342),
    .SET_B(net477),
    .Q(net498),
    .Q_N(net497));
 sky130_fd_sc_hd__mux4_4 c616 (.A0(net485),
    .A1(net975),
    .A2(clknet_1_0__leaf_net396),
    .A3(clknet_1_1__leaf_net394),
    .S0(net160),
    .S1(clknet_1_0__leaf_net881),
    .X(net499));
 sky130_fd_sc_hd__a221o_1 c617 (.A1(net451),
    .A2(net431),
    .B1(net420),
    .B2(net985),
    .C1(net1004),
    .X(net500));
 sky130_fd_sc_hd__sdfbbn_1 c618 (.CLK_N(clknet_4_10_0_clk),
    .D(net498),
    .RESET_B(clknet_1_0__leaf_net394),
    .SCD(net485),
    .SCE(net431),
    .SET_B(clknet_1_0__leaf_net739),
    .Q(net926));
 sky130_fd_sc_hd__mux4_2 c619 (.A0(net161),
    .A1(net471),
    .A2(clknet_1_1__leaf_net396),
    .A3(net284),
    .S0(net484),
    .S1(net951),
    .X(net501));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net3),
    .A1(net841),
    .A2(net862),
    .A3(net847),
    .S0(net863),
    .S1(net864),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net26),
    .A1(net832),
    .A2(net477),
    .A3(net946),
    .S0(clknet_1_1__leaf_net401),
    .S1(net671),
    .X(net880));
 sky130_fd_sc_hd__mux4_4 c621 (.A0(clknet_1_1__leaf_net329),
    .A1(net902),
    .A2(net164),
    .A3(net477),
    .S0(net935),
    .S1(net878),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net471),
    .A1(net903),
    .A2(net876),
    .A3(net884),
    .S0(net902),
    .S1(clknet_1_1__leaf_net493),
    .X(net503));
 sky130_fd_sc_hd__mux4_4 c623 (.A0(net501),
    .A1(clknet_1_1__leaf_net404),
    .A2(clknet_1_1__leaf_net394),
    .A3(net160),
    .S0(net973),
    .S1(net769),
    .X(net504));
 sky130_fd_sc_hd__mux4_2 c624 (.A0(net477),
    .A1(net284),
    .A2(net26),
    .A3(net451),
    .S0(net484),
    .S1(clknet_1_1__leaf_net739),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net431),
    .A1(net491),
    .A2(clknet_1_1__leaf_net329),
    .A3(net874),
    .S0(net164),
    .S1(net893),
    .X(net506));
 sky130_fd_sc_hd__mux4_2 c626 (.A0(net498),
    .A1(net26),
    .A2(net477),
    .A3(net284),
    .S0(clknet_1_1__leaf_net234),
    .S1(net764),
    .X(net507));
 sky130_fd_sc_hd__mux4_4 c627 (.A0(net893),
    .A1(net209),
    .A2(net875),
    .A3(clknet_1_1__leaf_net704),
    .S0(net771),
    .S1(net772),
    .X(net508));
 sky130_fd_sc_hd__mux4_2 c628 (.A0(net154),
    .A1(net884),
    .A2(net874),
    .A3(net26),
    .S0(clknet_1_1__leaf_net508),
    .S1(clknet_1_1__leaf_net757),
    .X(net509));
 sky130_fd_sc_hd__a221o_2 c629 (.A1(net377),
    .A2(clknet_1_1__leaf_net234),
    .B1(clknet_1_1__leaf_net394),
    .B2(net491),
    .C1(net772),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c63 (.A0(net863),
    .A1(net855),
    .A2(net829),
    .A3(net857),
    .S0(net864),
    .S1(net867),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c630 (.A0(clknet_1_1__leaf_net234),
    .A1(net893),
    .A2(clknet_1_0__leaf_net493),
    .A3(net930),
    .S0(clknet_1_0__leaf_net394),
    .S1(net933),
    .X(net511));
 sky130_fd_sc_hd__mux4_2 c631 (.A0(net946),
    .A1(clknet_1_0__leaf_net404),
    .A2(net714),
    .A3(net732),
    .S0(clknet_1_0__leaf_net739),
    .S1(net769),
    .X(net512));
 sky130_fd_sc_hd__sdfbbn_1 c632 (.CLK_N(clknet_4_9_0_clk),
    .D(net252),
    .RESET_B(net451),
    .SCD(net682),
    .SCE(clknet_1_0__leaf_net739),
    .SET_B(net769),
    .Q(net514),
    .Q_N(net513));
 sky130_fd_sc_hd__mux4_4 c633 (.A0(net507),
    .A1(clknet_1_1__leaf_net493),
    .A2(clknet_1_1__leaf_net508),
    .A3(clknet_1_1__leaf_net330),
    .S0(net715),
    .S1(net770),
    .X(net515));
 sky130_fd_sc_hd__mux4_2 c634 (.A0(clknet_1_1__leaf_net432),
    .A1(net873),
    .A2(net286),
    .A3(net513),
    .S0(clknet_1_0__leaf_net396),
    .S1(net769),
    .X(net516));
 sky130_fd_sc_hd__mux4_2 c635 (.A0(net252),
    .A1(net286),
    .A2(net514),
    .A3(clknet_1_1__leaf_net508),
    .S0(net672),
    .S1(net714),
    .X(net517));
 sky130_fd_sc_hd__a221oi_4 c636 (.A1(net451),
    .A2(net497),
    .B1(net161),
    .B2(clknet_1_1__leaf_net234),
    .C1(net772),
    .Y(net518));
 sky130_fd_sc_hd__mux4_2 c637 (.A0(net284),
    .A1(clknet_1_1__leaf_net234),
    .A2(net726),
    .A3(net769),
    .S0(net774),
    .S1(clknet_1_1__leaf_net775),
    .X(net871));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net850),
    .A1(net1),
    .A2(net867),
    .A3(net863),
    .S0(net859),
    .S1(net857),
    .X(net2));
 sky130_fd_sc_hd__or3b_1 c65 (.A(net833),
    .B(net811),
    .C_N(net817),
    .X(net3));
 sky130_fd_sc_hd__nor2_2 c66 (.A(net857),
    .B(net832),
    .Y(net4));
 sky130_fd_sc_hd__buf_6 c660 (.A(net733),
    .X(net519));
 sky130_fd_sc_hd__nor2b_1 c661 (.A(net198),
    .B_N(net70),
    .Y(net520));
 sky130_fd_sc_hd__clkinv_4 c662 (.A(net733),
    .Y(net521));
 sky130_fd_sc_hd__or2_1 c663 (.A(net947),
    .B(net521),
    .X(net522));
 sky130_fd_sc_hd__nor2_4 c664 (.A(net407),
    .B(net521),
    .Y(net523));
 sky130_fd_sc_hd__or2b_2 c665 (.A(net519),
    .B_N(net522),
    .X(net524));
 sky130_fd_sc_hd__or2_2 c666 (.A(net519),
    .B(net521),
    .X(net525));
 sky130_fd_sc_hd__or2b_4 c667 (.A(net524),
    .B_N(net410),
    .X(net526));
 sky130_fd_sc_hd__nand2_1 c668 (.A(net417),
    .B(net523),
    .Y(net527));
 sky130_fd_sc_hd__mux4_2 c669 (.A0(net526),
    .A1(net520),
    .A2(net521),
    .A3(net524),
    .S0(net519),
    .S1(net417),
    .X(net528));
 sky130_fd_sc_hd__nand2b_2 c67 (.A_N(net825),
    .B(net859),
    .Y(net889));
 sky130_fd_sc_hd__or2_1 c670 (.A(net524),
    .B(net762),
    .X(net529));
 sky130_fd_sc_hd__and2_1 c671 (.A(net529),
    .B(net525),
    .X(net530));
 sky130_fd_sc_hd__sdfbbp_1 c672 (.CLK(clknet_4_1_0_clk),
    .D(net529),
    .RESET_B(net519),
    .SCD(net521),
    .SCE(net527),
    .SET_B(net297),
    .Q(net532),
    .Q_N(net531));
 sky130_fd_sc_hd__buf_6 c673 (.A(net723),
    .X(net533));
 sky130_fd_sc_hd__a211oi_1 c674 (.A1(net522),
    .A2(net527),
    .B1(net298),
    .C1(net950),
    .Y(net534));
 sky130_fd_sc_hd__sdfbbn_1 c675 (.CLK_N(clknet_4_0_0_clk),
    .D(net297),
    .RESET_B(net532),
    .SCD(net525),
    .SCE(net421),
    .SET_B(net528),
    .Q(net536),
    .Q_N(net535));
 sky130_fd_sc_hd__inv_6 c676 (.A(net723),
    .Y(net537));
 sky130_fd_sc_hd__nand2b_4 c677 (.A_N(net520),
    .B(net950),
    .Y(net538));
 sky130_fd_sc_hd__a221o_1 c678 (.A1(net537),
    .A2(net538),
    .B1(net527),
    .C1(net762),
    .X(net539));
 sky130_fd_sc_hd__and2b_1 c679 (.A_N(net538),
    .B(net686),
    .X(net540));
 sky130_fd_sc_hd__nor2_1 c68 (.A(net945),
    .B(net855),
    .Y(net5));
 sky130_fd_sc_hd__sdfbbn_1 c680 (.CLK_N(clknet_4_1_0_clk),
    .D(net528),
    .RESET_B(net540),
    .SCD(net298),
    .SCE(net538),
    .SET_B(net686),
    .Q(net542),
    .Q_N(net541));
 sky130_fd_sc_hd__mux4_2 c681 (.A0(net537),
    .A1(net533),
    .A2(net540),
    .A3(net538),
    .S0(net686),
    .S1(net761),
    .X(net543));
 sky130_fd_sc_hd__a221oi_4 c682 (.A1(net531),
    .A2(net947),
    .B1(net523),
    .B2(net751),
    .C1(net765),
    .Y(net544));
 sky130_fd_sc_hd__a221oi_4 c683 (.A1(net540),
    .A2(net544),
    .B1(net87),
    .B2(net429),
    .C1(net535),
    .Y(net545));
 sky130_fd_sc_hd__a221o_2 c684 (.A1(net446),
    .A2(net817),
    .B1(net535),
    .B2(net531),
    .C1(net530),
    .X(net546));
 sky130_fd_sc_hd__a221oi_1 c685 (.A1(net536),
    .A2(clknet_1_0__leaf_net330),
    .B1(net521),
    .B2(net540),
    .C1(net525),
    .Y(net547));
 sky130_fd_sc_hd__sdfbbp_1 c686 (.CLK(clknet_4_0_0_clk),
    .D(net544),
    .RESET_B(net542),
    .SCD(clknet_1_0__leaf_net330),
    .SCE(net449),
    .SET_B(net546),
    .Q(net549),
    .Q_N(net548));
 sky130_fd_sc_hd__sdfbbn_1 c687 (.CLK_N(clknet_4_0_0_clk),
    .D(net991),
    .RESET_B(net524),
    .SCD(clknet_1_0__leaf_net447),
    .SCE(net530),
    .SET_B(net416),
    .Q(net551),
    .Q_N(net550));
 sky130_fd_sc_hd__sdfbbn_1 c688 (.CLK_N(clknet_4_1_0_clk),
    .D(net530),
    .RESET_B(net416),
    .SCD(net997),
    .SCE(net533),
    .SET_B(net538),
    .Q(net553),
    .Q_N(net552));
 sky130_fd_sc_hd__sdfbbp_1 c689 (.CLK(clknet_4_0_0_clk),
    .D(net410),
    .RESET_B(net546),
    .SCD(net446),
    .SCE(net541),
    .SET_B(net543),
    .Q(net555),
    .Q_N(net554));
 sky130_fd_sc_hd__nor2_2 c69 (.A(net829),
    .B(net857),
    .Y(net6));
 sky130_fd_sc_hd__mux4_2 c690 (.A0(net524),
    .A1(net555),
    .A2(net416),
    .A3(net550),
    .S0(net552),
    .S1(clknet_1_0__leaf_net330),
    .X(net556));
 sky130_fd_sc_hd__sdfbbn_1 c691 (.CLK_N(clknet_4_0_0_clk),
    .D(net996),
    .RESET_B(net410),
    .SCD(net543),
    .SCE(net416),
    .SET_B(clknet_1_0__leaf_net776),
    .Q(net558),
    .Q_N(net557));
 sky130_fd_sc_hd__mux4_2 c692 (.A0(clknet_1_1__leaf_net447),
    .A1(net947),
    .A2(net525),
    .A3(clknet_1_0__leaf_net219),
    .S0(clknet_1_0__leaf_net330),
    .S1(net530),
    .X(net559));
 sky130_fd_sc_hd__mux4_4 c693 (.A0(net532),
    .A1(net555),
    .A2(clknet_1_0__leaf_net330),
    .A3(net533),
    .S0(clknet_1_0__leaf_net776),
    .S1(clknet_1_0__leaf_net777),
    .X(net560));
 sky130_fd_sc_hd__a221o_1 c694 (.A1(net821),
    .A2(net410),
    .B1(net558),
    .B2(net554),
    .C1(net765),
    .X(net561));
 sky130_fd_sc_hd__sdfbbn_1 c695 (.CLK_N(clknet_4_0_0_clk),
    .D(net416),
    .RESET_B(net543),
    .SCD(net554),
    .SCE(net557),
    .SET_B(net987),
    .Q(net563),
    .Q_N(net562));
 sky130_fd_sc_hd__a221oi_1 c696 (.A1(net298),
    .A2(net410),
    .B1(net554),
    .B2(net765),
    .C1(net779),
    .Y(net564));
 sky130_fd_sc_hd__a221o_2 c697 (.A1(net558),
    .A2(net562),
    .B1(net297),
    .B2(net679),
    .C1(net733),
    .X(net565));
 sky130_fd_sc_hd__a221oi_2 c698 (.A1(net563),
    .A2(net524),
    .B1(net523),
    .B2(net733),
    .C1(net779),
    .Y(net566));
 sky130_fd_sc_hd__a221o_1 c699 (.A1(net563),
    .A2(net410),
    .B1(net765),
    .B2(clknet_1_1__leaf_net776),
    .C1(clknet_1_1__leaf_net777),
    .X(net567));
 sky130_fd_sc_hd__and3_1 c70 (.A(net5),
    .B(net859),
    .C(net946),
    .X(net7));
 sky130_fd_sc_hd__mux4_2 c700 (.A0(net566),
    .A1(net549),
    .A2(net555),
    .A3(clknet_1_0__leaf_net567),
    .S0(net436),
    .S1(net778),
    .X(net568));
 sky130_fd_sc_hd__mux4_4 c701 (.A0(net561),
    .A1(net551),
    .A2(clknet_1_0__leaf_net447),
    .A3(clknet_1_0__leaf_net568),
    .S0(net521),
    .S1(clknet_1_0__leaf_net567),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net555),
    .A1(net566),
    .A2(clknet_1_0__leaf_net568),
    .A3(clknet_1_0__leaf_net567),
    .S0(net723),
    .S1(net747),
    .X(net570));
 sky130_fd_sc_hd__a221o_2 c703 (.A1(net526),
    .A2(net561),
    .B1(clknet_1_0__leaf_net567),
    .B2(net679),
    .C1(net723),
    .X(net571));
 sky130_fd_sc_hd__sdfbbp_1 c704 (.CLK(clknet_4_1_0_clk),
    .D(net312),
    .RESET_B(net950),
    .SCD(clknet_1_0__leaf_net571),
    .SCE(net832),
    .SET_B(net975),
    .Q(net573),
    .Q_N(net572));
 sky130_fd_sc_hd__a21boi_1 c705 (.A1(net932),
    .A2(net538),
    .B1_N(net464),
    .Y(net574));
 sky130_fd_sc_hd__sdfbbn_2 c706 (.CLK_N(clknet_4_2_0_clk),
    .D(net574),
    .RESET_B(clknet_1_0__leaf_net571),
    .SCD(net523),
    .SCE(net565),
    .SET_B(net545),
    .Q(net576),
    .Q_N(net575));
 sky130_fd_sc_hd__a221o_4 c707 (.A1(net465),
    .A2(clknet_1_1__leaf_net567),
    .B1(net548),
    .B2(net932),
    .C1(net575),
    .X(net577));
 sky130_fd_sc_hd__mux4_2 c708 (.A0(net538),
    .A1(net525),
    .A2(net543),
    .A3(net943),
    .S0(net429),
    .S1(net575),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net565),
    .A1(net463),
    .A2(net546),
    .A3(net572),
    .S0(net575),
    .S1(net751),
    .X(net579));
 sky130_fd_sc_hd__or2b_1 c71 (.A(net851),
    .B_N(net857),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net542),
    .A1(net565),
    .A2(net449),
    .A3(net538),
    .S0(clknet_1_0__leaf_net568),
    .S1(net575),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net578),
    .A1(net573),
    .A2(net576),
    .A3(net947),
    .S0(net429),
    .S1(net780),
    .X(net581));
 sky130_fd_sc_hd__sedfxtp_1 c712 (.CLK(clknet_4_2_0_clk),
    .D(net553),
    .DE(net312),
    .SCD(net546),
    .SCE(net575),
    .Q(net582));
 sky130_fd_sc_hd__a211oi_4 c713 (.A1(net942),
    .A2(clknet_1_0__leaf_net568),
    .B1(net578),
    .C1(net575),
    .Y(net583));
 sky130_fd_sc_hd__a221oi_2 c714 (.A1(net95),
    .A2(net523),
    .B1(net541),
    .B2(net430),
    .C1(net575),
    .Y(net584));
 sky130_fd_sc_hd__sdfbbn_1 c715 (.CLK_N(clknet_4_3_0_clk),
    .D(net437),
    .RESET_B(net577),
    .SCD(net576),
    .SCE(net582),
    .SET_B(net565),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 c716 (.A(net729),
    .X(net587));
 sky130_fd_sc_hd__sdfbbp_1 c717 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net358),
    .RESET_B(net581),
    .SCD(net587),
    .SCE(net576),
    .SET_B(net994),
    .Q(net589),
    .Q_N(net588));
 sky130_fd_sc_hd__mux4_2 c718 (.A0(net525),
    .A1(net589),
    .A2(net545),
    .A3(net543),
    .S0(net553),
    .S1(clknet_1_0__leaf_net567),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net587),
    .A1(net589),
    .A2(net525),
    .A3(net575),
    .S0(net463),
    .S1(net546),
    .X(net591));
 sky130_fd_sc_hd__or2b_4 c72 (.A(net7),
    .B_N(net867),
    .X(net9));
 sky130_fd_sc_hd__mux4_4 c720 (.A0(net584),
    .A1(net586),
    .A2(net581),
    .A3(net589),
    .S0(net463),
    .S1(net526),
    .X(net592));
 sky130_fd_sc_hd__inv_1 c721 (.A(net729),
    .Y(net593));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net430),
    .A1(net589),
    .A2(net943),
    .A3(net575),
    .S0(net722),
    .S1(net783),
    .X(net594));
 sky130_fd_sc_hd__mux4_4 c723 (.A0(net449),
    .A1(net593),
    .A2(net594),
    .A3(net430),
    .S0(clknet_1_0__leaf_net330),
    .S1(net546),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net586),
    .A1(clknet_1_0__leaf_net219),
    .A2(net588),
    .A3(net575),
    .S0(net722),
    .S1(net751),
    .X(net596));
 sky130_fd_sc_hd__mux4_2 c725 (.A0(net549),
    .A1(net584),
    .A2(net588),
    .A3(net587),
    .S0(net785),
    .S1(net786),
    .X(net597));
 sky130_fd_sc_hd__mux4_4 c726 (.A0(clknet_1_1__leaf_net492),
    .A1(net207),
    .A2(clknet_1_1__leaf_net567),
    .A3(net933),
    .S0(net951),
    .S1(net768),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net87),
    .A1(net586),
    .A2(net943),
    .A3(net463),
    .S0(net130),
    .S1(net781),
    .X(net599));
 sky130_fd_sc_hd__mux4_2 c728 (.A0(net555),
    .A1(net594),
    .A2(net45),
    .A3(net526),
    .S0(net597),
    .S1(net491),
    .X(net600));
 sky130_fd_sc_hd__mux4_2 c729 (.A0(clknet_1_0__leaf_net590),
    .A1(net946),
    .A2(net576),
    .A3(net868),
    .S0(net782),
    .S1(net784),
    .X(net601));
 sky130_fd_sc_hd__and2_1 c73 (.A(net6),
    .B(net818),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net968),
    .A1(net302),
    .A2(net600),
    .A3(net932),
    .S0(net782),
    .S1(net786),
    .X(net602));
 sky130_fd_sc_hd__mux4_2 c731 (.A0(clknet_1_0__leaf_net370),
    .A1(net856),
    .A2(net130),
    .A3(net938),
    .S0(net302),
    .S1(net526),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net302),
    .A1(net582),
    .A2(net497),
    .A3(net600),
    .S0(net938),
    .S1(net998),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net472),
    .A1(clknet_1_0__leaf_net370),
    .A2(net523),
    .A3(net555),
    .S0(clknet_1_1__leaf_net330),
    .S1(net787),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_1__leaf_net567),
    .A1(net932),
    .A2(net378),
    .A3(net943),
    .S0(net576),
    .S1(net463),
    .X(net606));
 sky130_fd_sc_hd__mux4_2 c735 (.A0(net543),
    .A1(clknet_1_0__leaf_net370),
    .A2(net526),
    .A3(net600),
    .S0(net933),
    .S1(net789),
    .X(net607));
 sky130_fd_sc_hd__mux4_2 c736 (.A0(clknet_1_0__leaf_net489),
    .A1(net943),
    .A2(net526),
    .A3(net585),
    .S0(net788),
    .S1(net790),
    .X(net608));
 sky130_fd_sc_hd__sdfbbn_1 c737 (.CLK_N(clknet_4_8_0_clk),
    .D(clknet_1_0__leaf_net370),
    .RESET_B(net600),
    .SCD(clknet_1_1__leaf_net492),
    .SCE(net731),
    .SET_B(net790),
    .Q(net609));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(clknet_1_0__leaf_net608),
    .A1(clknet_1_1__leaf_net571),
    .A2(net523),
    .A3(net472),
    .S0(net554),
    .S1(net790),
    .X(net610));
 sky130_fd_sc_hd__mux4_2 c739 (.A0(net45),
    .A1(net968),
    .A2(net702),
    .A3(net768),
    .S0(net789),
    .S1(net791),
    .X(net611));
 sky130_fd_sc_hd__nor2_1 c74 (.A(net859),
    .B(net818),
    .Y(net11));
 sky130_fd_sc_hd__mux4_4 c740 (.A0(net609),
    .A1(net946),
    .A2(net611),
    .A3(net491),
    .S0(net933),
    .S1(net781),
    .X(net612));
 sky130_fd_sc_hd__mux4_2 c741 (.A0(net463),
    .A1(net472),
    .A2(net611),
    .A3(clknet_1_0__leaf_net492),
    .S0(net932),
    .S1(net725),
    .X(net613));
 sky130_fd_sc_hd__mux4_4 c742 (.A0(net597),
    .A1(net378),
    .A2(net611),
    .A3(net943),
    .S0(net731),
    .S1(net789),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net378),
    .A1(net612),
    .A2(net611),
    .A3(net463),
    .S0(clknet_1_1__leaf_net608),
    .S1(clknet_1_1__leaf_net590),
    .X(net615));
 sky130_fd_sc_hd__mux4_4 c744 (.A0(net856),
    .A1(clknet_1_1__leaf_net567),
    .A2(net600),
    .A3(net783),
    .S0(net784),
    .S1(net790),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net943),
    .A1(net543),
    .A2(clknet_1_1__leaf_net567),
    .A3(net611),
    .S0(net793),
    .S1(net794),
    .X(net617));
 sky130_fd_sc_hd__mux4_4 c746 (.A0(net130),
    .A1(net611),
    .A2(clknet_1_1__leaf_net567),
    .A3(net702),
    .S0(net793),
    .S1(net794),
    .X(net618));
 sky130_fd_sc_hd__mux4_2 c747 (.A0(net938),
    .A1(net617),
    .A2(net618),
    .A3(net378),
    .S0(clknet_1_0__leaf_net492),
    .S1(net786),
    .X(net619));
 sky130_fd_sc_hd__mux4_2 c748 (.A0(clknet_1_1__leaf_net568),
    .A1(net614),
    .A2(net164),
    .A3(net513),
    .S0(clknet_1_0__leaf_net493),
    .S1(net768),
    .X(net620));
 sky130_fd_sc_hd__mux4_4 c749 (.A0(net523),
    .A1(clknet_1_0__leaf_net493),
    .A2(net576),
    .A3(net600),
    .S0(net933),
    .S1(clknet_1_0__leaf_net508),
    .X(net621));
 sky130_fd_sc_hd__and3_2 c75 (.A(net811),
    .B(net861),
    .C(net832),
    .X(net12));
 sky130_fd_sc_hd__mux4_4 c750 (.A0(net491),
    .A1(net817),
    .A2(net576),
    .A3(net773),
    .S0(net792),
    .S1(clknet_1_0__leaf_net795),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(clknet_1_0__leaf_net508),
    .A1(clknet_1_0__leaf_net401),
    .A2(net526),
    .A3(clknet_1_0__leaf_net394),
    .S0(clknet_1_1__leaf_net795),
    .S1(clknet_1_0__leaf_net796),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net600),
    .A1(net576),
    .A2(clknet_1_0__leaf_net493),
    .A3(net207),
    .S0(clknet_1_0__leaf_net396),
    .S1(clknet_1_0__leaf_net796),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net514),
    .A1(clknet_1_0__leaf_net508),
    .A2(net286),
    .A3(clknet_1_1__leaf_net568),
    .S0(net676),
    .S1(net768),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net933),
    .A1(net576),
    .A2(net514),
    .A3(clknet_1_1__leaf_net330),
    .S0(clknet_1_0__leaf_net797),
    .S1(net798),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net526),
    .A1(net946),
    .A2(net773),
    .A3(clknet_1_0__leaf_net796),
    .S0(clknet_1_1__leaf_net797),
    .S1(net800),
    .X(net627));
 sky130_fd_sc_hd__mux4_4 c756 (.A0(clknet_1_0__leaf_net394),
    .A1(net498),
    .A2(net946),
    .A3(clknet_1_0__leaf_net508),
    .S0(clknet_1_0__leaf_net796),
    .S1(clknet_1_1__leaf_net797),
    .X(net628));
 sky130_fd_sc_hd__mux4_2 c757 (.A0(net627),
    .A1(clknet_1_0__leaf_net396),
    .A2(net286),
    .A3(net523),
    .S0(net933),
    .S1(clknet_1_0__leaf_net796),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net622),
    .A1(clknet_1_1__leaf_net330),
    .A2(net576),
    .A3(clknet_1_1__leaf_net796),
    .S0(clknet_1_0__leaf_net797),
    .S1(net800),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net946),
    .A1(clknet_1_1__leaf_net330),
    .A2(clknet_1_1__leaf_net568),
    .A3(net774),
    .S0(clknet_1_0__leaf_net775),
    .S1(net799),
    .X(net631));
 sky130_fd_sc_hd__nor2b_1 c76 (.A(net10),
    .B_N(net829),
    .Y(net13));
 sky130_fd_sc_hd__mux4_4 c760 (.A0(net286),
    .A1(clknet_1_0__leaf_net508),
    .A2(net732),
    .A3(net773),
    .S0(clknet_1_1__leaf_net797),
    .S1(net801),
    .X(net632));
 sky130_fd_sc_hd__mux4_4 c761 (.A0(net164),
    .A1(clknet_1_1__leaf_net493),
    .A2(clknet_1_0__leaf_net508),
    .A3(net676),
    .S0(net800),
    .S1(net802),
    .X(net633));
 sky130_fd_sc_hd__mux4_2 c762 (.A0(clknet_1_0__leaf_net704),
    .A1(net715),
    .A2(net724),
    .A3(clknet_1_0__leaf_net775),
    .S0(clknet_1_1__leaf_net796),
    .S1(net799));
 sky130_fd_sc_hd__and3_1 c77 (.A(net8),
    .B(net855),
    .C(net5),
    .X(net14));
 sky130_fd_sc_hd__a211o_1 c78 (.A1(net818),
    .A2(net11),
    .B1(net8),
    .C1(net823),
    .X(net15));
 sky130_fd_sc_hd__a211o_1 c79 (.A1(net14),
    .A2(net13),
    .B1(net4),
    .C1(net9),
    .X(net16));
 sky130_fd_sc_hd__a211o_1 c80 (.A1(net827),
    .A2(net9),
    .B1(net15),
    .C1(net836),
    .X(net17));
 sky130_fd_sc_hd__and3b_4 c81 (.A_N(net13),
    .B(net15),
    .C(net16),
    .X(net18));
 sky130_fd_sc_hd__nor2_1 c82 (.A(net9),
    .B(net13),
    .Y(net19));
 sky130_fd_sc_hd__a211oi_4 c83 (.A1(net15),
    .A2(net2),
    .B1(net9),
    .C1(net18),
    .Y(net20));
 sky130_fd_sc_hd__mux4_2 c84 (.A0(net11),
    .A1(net18),
    .A2(net20),
    .A3(net847),
    .S0(net945),
    .S1(net8),
    .X(net916));
 sky130_fd_sc_hd__nand2b_2 c85 (.A_N(net16),
    .B(net20),
    .Y(net21));
 sky130_fd_sc_hd__mux4_2 c86 (.A0(net17),
    .A1(net19),
    .A2(net21),
    .A3(net916),
    .S0(net20),
    .S1(net945),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c87 (.A0(net7),
    .A1(net21),
    .A2(net20),
    .A3(net17),
    .S0(net945),
    .S1(net916),
    .X(net23));
 sky130_fd_sc_hd__nor2b_4 c88 (.A(net867),
    .B_N(net823),
    .Y(net24));
 sky130_fd_sc_hd__nor2b_4 c89 (.A(net22),
    .B_N(net826),
    .Y(net25));
 sky130_fd_sc_hd__and2_4 c90 (.A(net14),
    .B(net18),
    .X(net26));
 sky130_fd_sc_hd__nand2b_1 c91 (.A_N(net26),
    .B(net25),
    .Y(net27));
 sky130_fd_sc_hd__nor3_1 c92 (.A(net836),
    .B(net27),
    .C(net867),
    .Y(net28));
 sky130_fd_sc_hd__nand2_1 c93 (.A(net45),
    .B(net22),
    .Y(net29));
 sky130_fd_sc_hd__nor2_1 c94 (.A(net866),
    .B(net946),
    .Y(net30));
 sky130_fd_sc_hd__and2b_1 c95 (.A_N(net27),
    .B(net30),
    .X(net31));
 sky130_fd_sc_hd__nor3_1 c96 (.A(net822),
    .B(net31),
    .C(net945),
    .Y(net32));
 sky130_fd_sc_hd__nor2_2 c97 (.A(net824),
    .B(net26),
    .Y(net33));
 sky130_fd_sc_hd__or3b_1 c98 (.A(net31),
    .B(net32),
    .C_N(net24),
    .X(net34));
 sky130_fd_sc_hd__nand2b_4 c99 (.A_N(net30),
    .B(net22),
    .Y(net35));
 sky130_fd_sc_hd__mux4_1 merge763 (.A0(net376),
    .A1(net458),
    .A2(clknet_1_1__leaf_net456),
    .A3(net481),
    .S0(clknet_1_1__leaf_net432),
    .S1(clknet_1_0__leaf_net881),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 merge764 (.A0(net199),
    .A1(net196),
    .A2(clknet_1_1__leaf_net219),
    .A3(net314),
    .S0(net298),
    .S1(net750),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_1 merge765 (.A(net727),
    .X(net636));
 sky130_fd_sc_hd__mux4_4 merge766 (.A0(net56),
    .A1(net925),
    .A2(net895),
    .A3(net165),
    .S0(net149),
    .S1(net692),
    .X(net637));
 sky130_fd_sc_hd__a221oi_1 merge767 (.A1(net205),
    .A2(net203),
    .B1(net85),
    .B2(net190),
    .C1(net938),
    .Y(net638));
 sky130_fd_sc_hd__a211o_1 merge768 (.A1(net845),
    .A2(net883),
    .B1(net109),
    .C1(net956),
    .X(net639));
 sky130_fd_sc_hd__a211oi_4 merge769 (.A1(net190),
    .A2(net297),
    .B1(clknet_1_0__leaf_net218),
    .C1(net214),
    .Y(net640));
 sky130_fd_sc_hd__a221oi_1 merge770 (.A1(net28),
    .A2(net145),
    .B1(net834),
    .B2(net892),
    .C1(net146),
    .Y(net641));
 sky130_fd_sc_hd__a211oi_1 merge771 (.A1(net298),
    .A2(net421),
    .B1(net416),
    .C1(net747),
    .Y(net642));
 sky130_fd_sc_hd__sdfbbn_1 merge772 (.CLK_N(clknet_4_12_0_clk),
    .D(net139),
    .RESET_B(net346),
    .SCD(clknet_1_1__leaf_net217),
    .SCE(net876),
    .SET_B(clknet_1_0__leaf_net738),
    .Q(net644),
    .Q_N(net643));
 sky130_fd_sc_hd__buf_16 merge773 (.A(net917),
    .X(net645));
 sky130_fd_sc_hd__mux4_1 merge774 (.A0(net248),
    .A1(net940),
    .A2(clknet_1_0__leaf_net254),
    .A3(net899),
    .S0(net252),
    .S1(net698),
    .X(net646));
 sky130_fd_sc_hd__a211oi_1 merge775 (.A1(net202),
    .A2(clknet_1_1__leaf_net219),
    .B1(net106),
    .C1(net942),
    .Y(net647));
 sky130_fd_sc_hd__a211oi_1 merge776 (.A1(net300),
    .A2(net821),
    .B1(net413),
    .C1(net303),
    .Y(net648));
 sky130_fd_sc_hd__sdfbbp_1 merge777 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net454),
    .RESET_B(clknet_1_0__leaf_net342),
    .SCD(clknet_1_0__leaf_net358),
    .SCE(net950),
    .SET_B(net749),
    .Q(net650),
    .Q_N(net649));
 sky130_fd_sc_hd__mux4_2 merge778 (.A0(clknet_1_0__leaf_net219),
    .A1(net552),
    .A2(net585),
    .A3(net546),
    .S0(net588),
    .S1(net785),
    .X(net651));
 sky130_fd_sc_hd__a221oi_2 merge779 (.A1(net338),
    .A2(net337),
    .B1(net341),
    .B2(net312),
    .C1(net189),
    .Y(net652));
 sky130_fd_sc_hd__a221o_1 merge780 (.A1(net300),
    .A2(net292),
    .B1(net939),
    .B2(net293),
    .C1(net306),
    .X(net653));
 sky130_fd_sc_hd__a221oi_4 merge781 (.A1(net290),
    .A2(net302),
    .B1(net190),
    .B2(net214),
    .C1(clknet_1_0__leaf_net218),
    .Y(net654));
 sky130_fd_sc_hd__sdfbbn_1 merge782 (.CLK_N(clknet_4_13_0_clk),
    .D(net90),
    .RESET_B(net154),
    .SCD(net145),
    .SCE(net23),
    .SET_B(net919),
    .Q(net656),
    .Q_N(net655));
 sky130_fd_sc_hd__a221o_1 merge783 (.A1(net417),
    .A2(net298),
    .B1(net442),
    .B2(net428),
    .C1(clknet_1_0__leaf_net439),
    .X(net657));
 sky130_fd_sc_hd__mux4_2 merge784 (.A0(clknet_1_0__leaf_net479),
    .A1(clknet_1_1__leaf_net489),
    .A2(net882),
    .A3(net884),
    .S0(net717),
    .S1(net767),
    .X(net658));
 sky130_fd_sc_hd__mux4_2 merge785 (.A0(net452),
    .A1(net451),
    .A2(net431),
    .A3(net237),
    .S0(net940),
    .S1(clknet_1_0__leaf_net241),
    .X(net659));
 sky130_fd_sc_hd__mux4_1 merge786 (.A0(net98),
    .A1(net88),
    .A2(net203),
    .A3(clknet_1_1__leaf_net241),
    .S0(net236),
    .S1(clknet_1_1__leaf_net219),
    .X(net660));
 sky130_fd_sc_hd__mux4_1 merge787 (.A0(net129),
    .A1(net244),
    .A2(net260),
    .A3(net351),
    .S0(net376),
    .S1(net712),
    .X(net661));
 sky130_fd_sc_hd__mux4_2 merge788 (.A0(net23),
    .A1(net892),
    .A2(net150),
    .A3(clknet_1_0__leaf_net256),
    .S0(net6),
    .S1(net976),
    .X(net662));
 sky130_fd_sc_hd__a211o_1 merge789 (.A1(net533),
    .A2(net528),
    .B1(net527),
    .C1(net530),
    .X(net663));
 sky130_fd_sc_hd__a221o_1 merge790 (.A1(net300),
    .A2(net312),
    .B1(net72),
    .B2(net407),
    .C1(net1000),
    .X(net664));
 sky130_fd_sc_hd__buf_6 merge791 (.A(net917),
    .X(net665));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net1005),
    .A1(net145),
    .A2(net56),
    .A3(net55),
    .S0(net888),
    .S1(net986),
    .X(net666));
 sky130_fd_sc_hd__mux4_2 merge793 (.A0(net966),
    .A1(net373),
    .A2(net376),
    .A3(clknet_1_1__leaf_net344),
    .S0(clknet_1_1__leaf_net367),
    .S1(net365),
    .X(net667));
 sky130_fd_sc_hd__a221oi_1 merge794 (.A1(net49),
    .A2(net44),
    .B1(net845),
    .B2(net857),
    .C1(net849),
    .Y(net668));
 sky130_fd_sc_hd__dfrbp_1 merge795 (.CLK(clknet_4_4_0_clk),
    .D(net323),
    .RESET_B(net332),
    .Q(net670),
    .Q_N(net669));
 sky130_fd_sc_hd__dfrbp_1 merge796 (.CLK(clknet_4_9_0_clk),
    .D(net499),
    .RESET_B(net500),
    .Q(net672),
    .Q_N(net671));
 sky130_fd_sc_hd__dfrtn_1 merge797 (.CLK_N(clknet_4_15_0_clk),
    .D(net173),
    .RESET_B(net174),
    .Q(net913));
 sky130_fd_sc_hd__and2_1 merge798 (.A(net191),
    .B(net192),
    .X(net673));
 sky130_fd_sc_hd__dfrtp_1 merge799 (.CLK(clknet_4_3_0_clk),
    .D(net468),
    .RESET_B(net473),
    .Q(net674));
 sky130_fd_sc_hd__nor2_1 merge800 (.A(net583),
    .B(net595),
    .Y(net675));
 sky130_fd_sc_hd__dfrtp_1 merge801 (.CLK(clknet_4_10_0_clk),
    .D(net620),
    .RESET_B(net623),
    .Q(net676));
 sky130_fd_sc_hd__and2_4 merge802 (.A(net364),
    .B(net379),
    .X(net677));
 sky130_fd_sc_hd__or2_2 merge803 (.A(net435),
    .B(net443),
    .X(net678));
 sky130_fd_sc_hd__dfrtp_1 merge804 (.CLK(clknet_4_0_0_clk),
    .D(net570),
    .RESET_B(net547),
    .Q(net679));
 sky130_fd_sc_hd__dfsbp_1 merge805 (.CLK(clknet_4_6_0_clk),
    .D(net339),
    .SET_B(net359),
    .Q(net681),
    .Q_N(net680));
 sky130_fd_sc_hd__dfsbp_1 merge806 (.CLK(clknet_4_9_0_clk),
    .D(net389),
    .SET_B(net391),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__dfstp_1 merge807 (.CLK(clknet_4_14_0_clk),
    .SET_B(net288),
    .Q(net879));
 sky130_fd_sc_hd__and2_4 merge808 (.A(net221),
    .B(net638),
    .X(net684));
 sky130_fd_sc_hd__dfstp_4 merge809 (.CLK(clknet_4_13_0_clk),
    .SET_B(net43),
    .Q(net908));
 sky130_fd_sc_hd__nand2b_1 merge810 (.A_N(net122),
    .B(net639),
    .Y(net685));
 sky130_fd_sc_hd__dfstp_1 merge811 (.CLK(clknet_4_1_0_clk),
    .D(net534),
    .Q(net539));
 sky130_fd_sc_hd__dlrbn_1 merge812 (.D(net159),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net155),
    .Q(net921),
    .Q_N(net687));
 sky130_fd_sc_hd__dlrbn_1 merge813 (.D(net653),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net301),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dlrbp_1 merge814 (.D(net647),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net243),
    .Q(net691),
    .Q_N(net690));
 sky130_fd_sc_hd__dlrbp_2 merge815 (.D(net668),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net57),
    .Q(net917),
    .Q_N(net692));
 sky130_fd_sc_hd__nor2_1 merge816 (.A(net598),
    .B(net599),
    .Y(net693));
 sky130_fd_sc_hd__dlrtn_2 merge817 (.D(net648),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net657),
    .Q(net694));
 sky130_fd_sc_hd__dlrtn_1 merge818 (.GATE_N(clknet_4_3_0_clk),
    .RESET_B(net486),
    .Q(net494));
 sky130_fd_sc_hd__dlrtn_1 merge819 (.D(net131),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net137));
 sky130_fd_sc_hd__dlrtp_1 merge820 (.D(net278),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net283),
    .Q(net697));
 sky130_fd_sc_hd__dlrtp_1 merge821 (.D(net249),
    .GATE(clknet_4_13_0_clk),
    .Q(net253));
 sky130_fd_sc_hd__dlrtp_1 merge822 (.D(net181),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net177),
    .Q(net909));
 sky130_fd_sc_hd__edfxbp_1 merge823 (.CLK(clknet_4_7_0_clk),
    .DE(net685),
    .Q(net700),
    .Q_N(net123));
 sky130_fd_sc_hd__and2b_2 merge824 (.A_N(net445),
    .B(net448),
    .X(net701));
 sky130_fd_sc_hd__edfxtp_1 merge825 (.CLK(clknet_4_8_0_clk),
    .D(net606),
    .DE(net607),
    .Q(net702));
 sky130_fd_sc_hd__or2b_1 merge826 (.A(net660),
    .B_N(net255),
    .X(net703));
 sky130_fd_sc_hd__sdlclkp_1 merge827 (.CLK(clknet_4_11_0_clk),
    .GATE(net506),
    .SCE(net633),
    .GCLK(net704));
 sky130_fd_sc_hd__or2_4 merge828 (.A(net393),
    .B(net518),
    .X(net705));
 sky130_fd_sc_hd__sdlclkp_2 merge829 (.CLK(clknet_4_7_0_clk),
    .GATE(net223),
    .SCE(net684),
    .GCLK(net706));
 sky130_fd_sc_hd__sdlclkp_4 merge830 (.CLK(clknet_4_5_0_clk),
    .GATE(net333),
    .SCE(net640),
    .GCLK(net707));
 sky130_fd_sc_hd__dfrbp_1 merge831 (.CLK(clknet_4_13_0_clk),
    .D(net661),
    .RESET_B(net666),
    .Q(net709),
    .Q_N(net708));
 sky130_fd_sc_hd__dfrbp_1 merge832 (.CLK(clknet_4_4_0_clk),
    .D(net678),
    .RESET_B(net635),
    .Q(net711),
    .Q_N(net710));
 sky130_fd_sc_hd__dfrtn_1 merge833 (.CLK_N(clknet_4_12_0_clk),
    .D(net677),
    .RESET_B(net652),
    .Q(net712));
 sky130_fd_sc_hd__dfrtp_4 merge834 (.CLK(clknet_4_5_0_clk),
    .D(net703),
    .RESET_B(net673),
    .Q(net713));
 sky130_fd_sc_hd__dfrtp_1 merge835 (.CLK(clknet_4_9_0_clk),
    .D(net509),
    .RESET_B(net516),
    .Q(net714));
 sky130_fd_sc_hd__dfrtp_1 merge836 (.CLK(clknet_4_11_0_clk),
    .D(net510),
    .RESET_B(net632),
    .Q(net715));
 sky130_fd_sc_hd__dfsbp_1 merge837 (.CLK(clknet_4_9_0_clk),
    .D(net262),
    .SET_B(net360),
    .Q(net717),
    .Q_N(net716));
 sky130_fd_sc_hd__and2_2 merge838 (.A(net179),
    .B(net397),
    .X(net718));
 sky130_fd_sc_hd__dfsbp_1 merge839 (.CLK(clknet_4_7_0_clk),
    .D(net654),
    .SET_B(net345),
    .Q(net720),
    .Q_N(net719));
 sky130_fd_sc_hd__dfstp_1 merge840 (.CLK(clknet_4_15_0_clk),
    .D(net178),
    .SET_B(net162),
    .Q(net721));
 sky130_fd_sc_hd__dfstp_2 merge841 (.CLK(clknet_4_1_0_clk),
    .D(net675),
    .SET_B(net664),
    .Q(net722));
 sky130_fd_sc_hd__dfstp_2 merge842 (.CLK(clknet_4_0_0_clk),
    .D(net663),
    .SET_B(net569),
    .Q(net723));
 sky130_fd_sc_hd__dlrbn_1 merge843 (.D(net601),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net631),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__dlrbn_1 merge844 (.D(net400),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net705),
    .Q(net890),
    .Q_N(net726));
 sky130_fd_sc_hd__dlrbp_1 merge845 (.D(net641),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net662),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__dlrbp_1 merge846 (.D(net701),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net651),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dlrtn_1 merge847 (.D(net602),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net693),
    .Q(net731));
 sky130_fd_sc_hd__dlrtn_1 merge848 (.D(net629),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net511),
    .Q(net732));
 sky130_fd_sc_hd__dlrtn_2 merge849 (.D(net564),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net642),
    .Q(net733));
 sky130_fd_sc_hd__dlrtp_2 merge850 (.D(net168),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net718),
    .Q(net734));
 sky130_fd_sc_hd__dfxbp_1 s851 (.CLK(clknet_4_13_0_clk),
    .D(net141),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__dfxbp_1 s852 (.CLK(clknet_4_14_0_clk),
    .D(net143),
    .Q(net894),
    .Q_N(net737));
 sky130_fd_sc_hd__dfxtp_2 s853 (.CLK(clknet_4_15_0_clk),
    .D(net152),
    .Q(net919));
 sky130_fd_sc_hd__dfxtp_2 s854 (.CLK(clknet_4_15_0_clk),
    .D(net169),
    .Q(net896));
 sky130_fd_sc_hd__dfxtp_1 s855 (.CLK(clknet_4_14_0_clk),
    .D(net180),
    .Q(net924));
 sky130_fd_sc_hd__dlclkp_1 s856 (.CLK(clknet_4_12_0_clk),
    .GATE(net246),
    .GCLK(net881));
 sky130_fd_sc_hd__dlclkp_2 s857 (.CLK(clknet_4_13_0_clk),
    .GATE(net265),
    .GCLK(net738));
 sky130_fd_sc_hd__dlclkp_4 s858 (.CLK(clknet_4_12_0_clk),
    .GATE(net272),
    .GCLK(net739));
 sky130_fd_sc_hd__dlxbn_1 s859 (.D(net277),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net741),
    .Q_N(net740));
 sky130_fd_sc_hd__dlxbn_1 s860 (.D(net279),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net743),
    .Q_N(net742));
 sky130_fd_sc_hd__dlxbp_1 s861 (.D(net281),
    .GATE(clknet_4_14_0_clk),
    .Q(net745),
    .Q_N(net744));
 sky130_fd_sc_hd__dlxtn_1 s862 (.D(net287),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net915));
 sky130_fd_sc_hd__dlxtn_2 s863 (.D(net310),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net746));
 sky130_fd_sc_hd__dlxtn_4 s864 (.D(net311),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net747));
 sky130_fd_sc_hd__dlxtp_1 s865 (.D(net322),
    .GATE(clknet_4_7_0_clk),
    .Q(net748));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s866 (.D(net334),
    .SLEEP_B(clknet_4_5_0_clk),
    .Q(net749));
 sky130_fd_sc_hd__dfxbp_2 s867 (.CLK(clknet_4_4_0_clk),
    .D(net335),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__dfxbp_1 s868 (.CLK(clknet_4_6_0_clk),
    .D(net353),
    .Q(net753),
    .Q_N(net752));
 sky130_fd_sc_hd__dfxtp_1 s869 (.CLK(clknet_4_6_0_clk),
    .D(net356),
    .Q(net754));
 sky130_fd_sc_hd__dfxtp_2 s870 (.CLK(clknet_4_9_0_clk),
    .D(net357),
    .Q(net755));
 sky130_fd_sc_hd__dfxtp_1 s871 (.CLK(clknet_4_12_0_clk),
    .D(net369),
    .Q(net756));
 sky130_fd_sc_hd__dlclkp_1 s872 (.CLK(clknet_4_9_0_clk),
    .GATE(net382),
    .GCLK(net757));
 sky130_fd_sc_hd__dlclkp_2 s873 (.CLK(clknet_4_9_0_clk),
    .GATE(net383),
    .GCLK(net758));
 sky130_fd_sc_hd__dlclkp_4 s874 (.CLK(clknet_4_14_0_clk),
    .GATE(net395),
    .GCLK(net886));
 sky130_fd_sc_hd__dlxbn_1 s875 (.D(net425),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net760),
    .Q_N(net759));
 sky130_fd_sc_hd__dlxbn_1 s876 (.D(net426),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net762),
    .Q_N(net761));
 sky130_fd_sc_hd__dlxbp_1 s877 (.D(net427),
    .GATE(clknet_4_4_0_clk),
    .Q(net764),
    .Q_N(net763));
 sky130_fd_sc_hd__dlxtn_2 s878 (.D(net440),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net765));
 sky130_fd_sc_hd__dlxtn_1 s879 (.D(net450),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net766));
 sky130_fd_sc_hd__dlxtn_1 s880 (.D(net475),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net767));
 sky130_fd_sc_hd__dlxtp_1 s881 (.D(net487),
    .GATE(clknet_4_8_0_clk),
    .Q(net768));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s882 (.D(net502),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net769));
 sky130_fd_sc_hd__dfxbp_1 s883 (.CLK(clknet_4_11_0_clk),
    .D(net503),
    .Q(net877));
 sky130_fd_sc_hd__dfxbp_1 s884 (.CLK(clknet_4_11_0_clk),
    .D(net504),
    .Q(net771),
    .Q_N(net770));
 sky130_fd_sc_hd__dfxtp_1 s885 (.CLK(clknet_4_11_0_clk),
    .D(net505),
    .Q(net772));
 sky130_fd_sc_hd__dfxtp_1 s886 (.CLK(clknet_4_11_0_clk),
    .D(net512),
    .Q(net773));
 sky130_fd_sc_hd__dfxtp_1 s887 (.CLK(clknet_4_11_0_clk),
    .D(net515),
    .Q(net774));
 sky130_fd_sc_hd__dlclkp_1 s888 (.CLK(clknet_4_11_0_clk),
    .GATE(net517),
    .GCLK(net775));
 sky130_fd_sc_hd__dlclkp_2 s889 (.CLK(clknet_4_0_0_clk),
    .GATE(net556),
    .GCLK(net776));
 sky130_fd_sc_hd__dlclkp_4 s890 (.CLK(clknet_4_0_0_clk),
    .GATE(net559),
    .GCLK(net777));
 sky130_fd_sc_hd__dlxbn_1 s891 (.D(net560),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net779),
    .Q_N(net778));
 sky130_fd_sc_hd__dlxbn_1 s892 (.D(net579),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dlxbp_1 s893 (.D(net580),
    .GATE(clknet_4_2_0_clk),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__dlxtn_1 s894 (.D(net591),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net784));
 sky130_fd_sc_hd__dlxtn_1 s895 (.D(net592),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net785));
 sky130_fd_sc_hd__dlxtn_1 s896 (.D(net596),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net786));
 sky130_fd_sc_hd__dlxtp_1 s897 (.D(net603),
    .GATE(clknet_4_2_0_clk),
    .Q(net787));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s898 (.D(net604),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net788));
 sky130_fd_sc_hd__dfxbp_1 s899 (.CLK(clknet_4_2_0_clk),
    .D(net605),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dfxbp_1 s900 (.CLK(clknet_4_2_0_clk),
    .D(net610),
    .Q(net791));
 sky130_fd_sc_hd__dfxtp_1 s901 (.CLK(clknet_4_8_0_clk),
    .D(net613),
    .Q(net792));
 sky130_fd_sc_hd__dfxtp_1 s902 (.CLK(clknet_4_2_0_clk),
    .D(net615),
    .Q(net793));
 sky130_fd_sc_hd__dfxtp_1 s903 (.CLK(clknet_4_2_0_clk),
    .D(net616),
    .Q(net794));
 sky130_fd_sc_hd__dlclkp_1 s904 (.CLK(clknet_4_10_0_clk),
    .GATE(net619),
    .GCLK(net795));
 sky130_fd_sc_hd__dlclkp_2 s905 (.CLK(clknet_4_8_0_clk),
    .GATE(net621),
    .GCLK(net796));
 sky130_fd_sc_hd__dlclkp_4 s906 (.CLK(clknet_4_10_0_clk),
    .GATE(net624),
    .GCLK(net797));
 sky130_fd_sc_hd__dlxbn_1 s907 (.D(net625),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net798));
 sky130_fd_sc_hd__dlxbn_1 s908 (.D(net626),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dlxbp_1 s909 (.D(net628),
    .GATE(clknet_4_10_0_clk),
    .Q(net801));
 sky130_fd_sc_hd__dlxtn_1 s910 (.D(net630),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net802));
 sky130_fd_sc_hd__dlxtn_1 s911 (.D(net634),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net803));
 sky130_fd_sc_hd__dlxtn_1 s912 (.D(net637),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net804));
 sky130_fd_sc_hd__dlxtp_1 s913 (.D(net646),
    .GATE(clknet_4_12_0_clk),
    .Q(net805));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s914 (.D(net658),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net806));
 sky130_fd_sc_hd__dfxbp_1 s915 (.CLK(clknet_4_6_0_clk),
    .D(net659),
    .Q(net808),
    .Q_N(net807));
 sky130_fd_sc_hd__dfxbp_1 s916 (.CLK(clknet_4_12_0_clk),
    .D(net667),
    .Q(net810),
    .Q_N(net809));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(in0),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net814));
 sky130_fd_sc_hd__buf_12 input7 (.A(in14),
    .X(net815));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net816));
 sky130_fd_sc_hd__buf_4 input9 (.A(in16),
    .X(net817));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in18),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net820));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net821));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net822));
 sky130_fd_sc_hd__buf_4 input15 (.A(in21),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in22),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in23),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in25),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in26),
    .X(net828));
 sky130_fd_sc_hd__buf_1 input21 (.A(in27),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(in28),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_8 input24 (.A(in3),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(in31),
    .X(net834));
 sky130_fd_sc_hd__buf_2 input27 (.A(in32),
    .X(net835));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net836));
 sky130_fd_sc_hd__buf_2 input29 (.A(in34),
    .X(net837));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(in36),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(in37),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in38),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in39),
    .X(net842));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(in4),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(in40),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(in41),
    .X(net845));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net846));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net847));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net849));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(in47),
    .X(net851));
 sky130_fd_sc_hd__buf_1 input44 (.A(in48),
    .X(net852));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(in5),
    .X(net854));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(in50),
    .X(net855));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net856));
 sky130_fd_sc_hd__buf_2 input49 (.A(in52),
    .X(net857));
 sky130_fd_sc_hd__buf_1 input50 (.A(in53),
    .X(net858));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(in54),
    .X(net859));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(in55),
    .X(net860));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(in57),
    .X(net862));
 sky130_fd_sc_hd__buf_1 input55 (.A(in58),
    .X(net863));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(in59),
    .X(net864));
 sky130_fd_sc_hd__buf_1 input57 (.A(in6),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(in60),
    .X(net866));
 sky130_fd_sc_hd__buf_4 input59 (.A(in61),
    .X(net867));
 sky130_fd_sc_hd__buf_4 input60 (.A(in7),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in8),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in9),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net871),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output64 (.A(net207),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net873),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net874),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output67 (.A(net875),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output68 (.A(net876),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net877),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net878),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net879),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net880),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(clknet_1_1__leaf_net881),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output74 (.A(net882),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net883),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output76 (.A(net884),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output77 (.A(net885),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(clknet_1_1__leaf_net886),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output79 (.A(net887),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net888),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output81 (.A(net889),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output82 (.A(net890),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output83 (.A(net891),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output84 (.A(net892),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output85 (.A(net893),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output86 (.A(net894),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output87 (.A(net895),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output88 (.A(net896),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output89 (.A(net897),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output90 (.A(net898),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output91 (.A(net899),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output92 (.A(net900),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output93 (.A(net901),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output94 (.A(net902),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output95 (.A(net903),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net904),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output97 (.A(net905),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net906),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output99 (.A(net950),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output100 (.A(net908),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output101 (.A(net909),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output102 (.A(net910),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output103 (.A(net911),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output104 (.A(net320),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output105 (.A(net913),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output106 (.A(net914),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output107 (.A(net915),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net916),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output109 (.A(net917),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output110 (.A(net918),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output111 (.A(net919),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output112 (.A(net920),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output113 (.A(net921),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output114 (.A(net922),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output115 (.A(net923),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output116 (.A(net924),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output117 (.A(net925),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output118 (.A(net926),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output119 (.A(net927),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output120 (.A(net928),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(net244),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_2 max_cap122 (.A(net928),
    .X(net930));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net138),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_2 max_cap124 (.A(net545),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(net885),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_2 max_cap126 (.A(net117),
    .X(net934));
 sky130_fd_sc_hd__buf_12 fanout127 (.A(net912),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net189),
    .X(net936));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net927),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(net84),
    .X(net938));
 sky130_fd_sc_hd__buf_12 fanout131 (.A(net80),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_8 fanout132 (.A(net235),
    .X(net940));
 sky130_fd_sc_hd__buf_1 max_cap133 (.A(net105),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_2 max_cap134 (.A(net70),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net349),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_2 max_cap136 (.A(net1003),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net889),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net4),
    .X(net946));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net194),
    .X(net947));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net949),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__buf_6 fanout142 (.A(net907),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_8 fanout143 (.A(net907),
    .X(net951));
 sky130_fd_sc_hd__buf_12 fanout144 (.A(net64),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 fanout145 (.A(net955),
    .X(net953));
 sky130_fd_sc_hd__buf_1 fanout146 (.A(net955),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net103),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_2 fanout149 (.A(net103),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_8 fanout150 (.A(net849),
    .X(net958));
 sky130_fd_sc_hd__inv_8 c291_1 (.A(clknet_1_0__leaf_net706),
    .Y(net959));
 sky130_fd_sc_hd__inv_8 net899_2 (.A(clknet_1_0__leaf_net706),
    .Y(net960));
 sky130_fd_sc_hd__inv_8 net899_3 (.A(clknet_1_0__leaf_net706),
    .Y(net961));
 sky130_fd_sc_hd__inv_1 c293_5 (.A(clknet_1_0__leaf_net706),
    .Y(net963));
 sky130_fd_sc_hd__inv_1 c293_6 (.A(clknet_1_0__leaf_net706),
    .Y(net964));
 sky130_fd_sc_hd__inv_1 c293_7 (.A(clknet_1_0__leaf_net706),
    .Y(net965));
 sky130_fd_sc_hd__inv_6 c425_9 (.A(clknet_1_1__leaf_net707),
    .Y(net967));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net797 (.A(net797),
    .X(clknet_0_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_0__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_1__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net796 (.A(net796),
    .X(clknet_0_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_0__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_1__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net795 (.A(net795),
    .X(clknet_0_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net795 (.A(clknet_0_net795),
    .X(clknet_1_0__leaf_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net795 (.A(clknet_0_net795),
    .X(clknet_1_1__leaf_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net777 (.A(net777),
    .X(clknet_0_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_0__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_1__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net567 (.A(net567),
    .X(clknet_0_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_0__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net590 (.A(net590),
    .X(clknet_0_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net590 (.A(clknet_0_net590),
    .X(clknet_1_0__leaf_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net590 (.A(clknet_0_net590),
    .X(clknet_1_1__leaf_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net571 (.A(net571),
    .X(clknet_0_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_0__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_1__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net568 (.A(net568),
    .X(clknet_0_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_0__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_1__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net776 (.A(net776),
    .X(clknet_0_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net776 (.A(clknet_0_net776),
    .X(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net776 (.A(clknet_0_net776),
    .X(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net775 (.A(net775),
    .X(clknet_0_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_0__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net886 (.A(net886),
    .X(clknet_0_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net886 (.A(clknet_0_net886),
    .X(clknet_1_0__leaf_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net886 (.A(clknet_0_net886),
    .X(clknet_1_1__leaf_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net401 (.A(net401),
    .X(clknet_0_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_0__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net758 (.A(net758),
    .X(clknet_0_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_0__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_1__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net608 (.A(net608),
    .X(clknet_0_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_0__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_1__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net493 (.A(net493),
    .X(clknet_0_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_0__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_1__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net704 (.A(net704),
    .X(clknet_0_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net704 (.A(clknet_0_net704),
    .X(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net704 (.A(clknet_0_net704),
    .X(clknet_1_1__leaf_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net508 (.A(net508),
    .X(clknet_0_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_0__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_1__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net492 (.A(net492),
    .X(clknet_0_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_0__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_1__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net488 (.A(net488),
    .X(clknet_0_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_0__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_1__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net757 (.A(net757),
    .X(clknet_0_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_0__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_1__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net739 (.A(net739),
    .X(clknet_0_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net739 (.A(clknet_0_net739),
    .X(clknet_1_0__leaf_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net739 (.A(clknet_0_net739),
    .X(clknet_1_1__leaf_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net738 (.A(net738),
    .X(clknet_0_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net738 (.A(clknet_0_net738),
    .X(clknet_1_0__leaf_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net738 (.A(clknet_0_net738),
    .X(clknet_1_1__leaf_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net266 (.A(net266),
    .X(clknet_0_net266));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net266 (.A(clknet_0_net266),
    .X(clknet_1_0__leaf_net266));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net266 (.A(clknet_0_net266),
    .X(clknet_1_1__leaf_net266));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net370 (.A(net370),
    .X(clknet_0_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_0__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net881 (.A(net881),
    .X(clknet_0_net881));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net881 (.A(clknet_0_net881),
    .X(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net881 (.A(clknet_0_net881),
    .X(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net707 (.A(net707),
    .X(clknet_0_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_0__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_1__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net331 (.A(net331),
    .X(clknet_0_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_0__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_1__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net706 (.A(net706),
    .X(clknet_0_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net247 (.A(net247),
    .X(clknet_0_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net217 (.A(net217),
    .X(clknet_0_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_1__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net439 (.A(net439),
    .X(clknet_0_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_0__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_1__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net394 (.A(net394),
    .X(clknet_0_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_0__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_1__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net329 (.A(net329),
    .X(clknet_0_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net447 (.A(net447),
    .X(clknet_0_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_0__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_1__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net432 (.A(net432),
    .X(clknet_0_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net432 (.A(clknet_0_net432),
    .X(clknet_1_0__leaf_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net432 (.A(clknet_0_net432),
    .X(clknet_1_1__leaf_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net358 (.A(net358),
    .X(clknet_0_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_0__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_1__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net344 (.A(net344),
    .X(clknet_0_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net344 (.A(clknet_0_net344),
    .X(clknet_1_0__leaf_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net344 (.A(clknet_0_net344),
    .X(clknet_1_1__leaf_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net330 (.A(net330),
    .X(clknet_0_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net240 (.A(net240),
    .X(clknet_0_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net240 (.A(clknet_0_net240),
    .X(clknet_1_0__leaf_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net240 (.A(clknet_0_net240),
    .X(clknet_1_1__leaf_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net342 (.A(net342),
    .X(clknet_0_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net241 (.A(net241),
    .X(clknet_0_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_1__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net219 (.A(net219),
    .X(clknet_0_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net256 (.A(net256),
    .X(clknet_0_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_0__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_1__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net218 (.A(net218),
    .X(clknet_0_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_1__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net234 (.A(net234),
    .X(clknet_0_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net232 (.A(net232),
    .X(clknet_0_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net454 (.A(net454),
    .X(clknet_0_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_0__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_1__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net456 (.A(net456),
    .X(clknet_0_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_0__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_1__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net239 (.A(net239),
    .X(clknet_0_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net239 (.A(clknet_0_net239),
    .X(clknet_1_0__leaf_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net239 (.A(clknet_0_net239),
    .X(clknet_1_1__leaf_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net254 (.A(net254),
    .X(clknet_0_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_0__leaf_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_1__leaf_net254));
 sky130_fd_sc_hd__and2b_4 clone1 (.A_N(net822),
    .B(net975),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net912),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net209),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net64),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1007),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net80),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net79),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net907),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_1 clone9 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net912),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_4 clone11 (.A(net64),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net939),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net976),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net976),
    .X(net978));
 sky130_fd_sc_hd__buf_2 rebuffer15 (.A(net204),
    .X(net979));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer16 (.A(net979),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net251),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net756),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net735),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net778),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net688),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net408),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net924),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net521),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net472),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net919),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net554),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net755),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net551),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net536),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net786),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net304),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net713),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net354),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net909),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net748),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net764),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net150),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net697),
    .X(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_C (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_Y (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_D (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SCE (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_SCD (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_D (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B_N (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_SET_B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_RESET_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_SCD (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_Y (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_Q_N (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_X (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_C1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_C1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_Y (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_Y (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SCD (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_DE (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_SCD (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_Y (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_SCE (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_X (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net234_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_Y (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_C_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_Y (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_C1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_Y (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_RESET_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_S0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_D (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_SCE (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_Q_N (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_Q (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_D (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_Y (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_X (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCE (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_X (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_C1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_C1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1_N (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Y (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_B1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_D (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SET_B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A3 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_Y (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_S0 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_SCD (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S0 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_C1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S0 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A3 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_X (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_B2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_DE (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_D (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_SCE (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_RESET_B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_SCE (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_RESET_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_Q_N (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_Y (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A_N (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net330_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_D (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_D (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_Q (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_D (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_C (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_Q (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_Y (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A_N (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold25_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_D (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_DE (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A2 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_Y (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SCE (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_SCD (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_RESET_B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_Y (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_RESET_B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_D (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B_N (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_SET_B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_B1_N (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_Q_N (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_B1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_D (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_SCE (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_RESET_B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_SET_B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_SCD (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_Y (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_B1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Q_N (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SCD (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_RESET_B (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_X (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_SCE (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SCD (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B1_N (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_Y (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_Q_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_D (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_Q (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A0 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_X (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_RESET_B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SCE (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SET_B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_RESET_B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_Y (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_SCD (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_RESET_B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_SET_B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_X (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_Q (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold28_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SET_B (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_Q (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_SET_B (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B2 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B1_N (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_Y (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B2 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_X (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_Q_N (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_C (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_Y (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_SCD (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_Y (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_C1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_SCD (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A0 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_SET_B (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A3 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_SCE (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A_N (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_Y (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_RESET_B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_SCD (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SET_B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_X (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SCD (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_B2 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_Q_N (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_Q (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_SCE (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCD (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_Q (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_Y (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_Y (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone11_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_D (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_C (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold36_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_Q (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_SET_B (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_C1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_Q (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_Q (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_C1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_C1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_C1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_C1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_Q (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_C1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_C1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_C1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_C1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_C1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_SET_B (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_D (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B1_N (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_Y (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_Y (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_C1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_D (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_SCD (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_Y (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_C1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_Y (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_C1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B_N (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_SCD (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_S (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_C_N (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_A_N (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A_N (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B_N (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_C1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A_N (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A_N (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B1_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_C (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_SCE (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1_N (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B_N (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_C (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_C (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SCE (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_B1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_D (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_B1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_C1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_B2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B_N (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A_N (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A_N (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_C (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B_N (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Q (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_SCE (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_C1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_Q (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCD (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SCD (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_C1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_Y (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_RESET_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_B2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_Y (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_B1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_C1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_Y (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_C1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_B1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_Y (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_B2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_B1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_Y (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_Y (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_Q (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B_N (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_Y (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_Q (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_C (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B_N (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_Q (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_C_N (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold29_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_Q (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_SET_B (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_B1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_C1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_Y (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap122_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_Y (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_RESET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_C1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_D (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_B1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap122_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_B1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B1_N (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_C1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_C (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_B1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_B1_N (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B1_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_C1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_C (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_C (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_C1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_C1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_B1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_C (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_B1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap134_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_C1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCE (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap136_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_B2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_C1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_B1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_C1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_C (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SCD (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_C (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_C1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B1_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_SCD (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_C1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_C_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_C1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B1_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_SCE (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_RESET_B (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_C1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_B2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_C1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_C (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_C (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_C1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_C (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_C1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_C1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_C (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_C1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B2 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SET_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A_N (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_SLEEP_B (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B2 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_B1_N (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_S1 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net881_X (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net881_X (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_C1 (.DIODE(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net217_X (.DIODE(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1_N (.DIODE(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net329_X (.DIODE(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net329_X (.DIODE(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net330_A (.DIODE(clknet_0_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net330_A (.DIODE(clknet_0_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net330_X (.DIODE(clknet_0_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_C1 (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SET_B (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_SCE (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_SCE (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCE (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A2 (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_SCD (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S1 (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net330_X (.DIODE(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SCD (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_SCE (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCE (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net330_X (.DIODE(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A0 (.DIODE(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net219_X (.DIODE(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_S0 (.DIODE(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A2 (.DIODE(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A2 (.DIODE(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S1 (.DIODE(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net219_X (.DIODE(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B1_N (.DIODE(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_C1 (.DIODE(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net234_X (.DIODE(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_B2 (.DIODE(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net234_X (.DIODE(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone9_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone9_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCD (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SET_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone11_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B_N (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_B2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_RESET_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold25_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net9));
 sky130_fd_sc_hd__and2b_1 clone2 (.A_N(net822),
    .B(net952),
    .X(net981));
 sky130_fd_sc_hd__and2b_1 clone3 (.A_N(net819),
    .B(net823),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_1 clone4 (.A(net64),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net200),
    .X(net1007));
 sky130_fd_sc_hd__a211o_1 clone10 (.A1(net854),
    .A2(net66),
    .B1(net868),
    .C1(net948),
    .X(net1008));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
