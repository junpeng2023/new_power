module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net631;
 wire clknet_1_0__leaf_net631;
 wire clknet_1_1__leaf_net631;
 wire clknet_0_net726;
 wire clknet_1_0__leaf_net726;
 wire clknet_1_1__leaf_net726;
 wire clknet_0_net708;
 wire clknet_1_0__leaf_net708;
 wire clknet_1_1__leaf_net708;
 wire clknet_0_net610;
 wire clknet_1_0__leaf_net610;
 wire clknet_1_1__leaf_net610;
 wire clknet_0_net707;
 wire clknet_1_0__leaf_net707;
 wire clknet_1_1__leaf_net707;
 wire clknet_0_net615;
 wire clknet_1_0__leaf_net615;
 wire clknet_1_1__leaf_net615;
 wire clknet_0_net592;
 wire clknet_1_0__leaf_net592;
 wire clknet_1_1__leaf_net592;
 wire clknet_0_net691;
 wire clknet_1_0__leaf_net691;
 wire clknet_1_1__leaf_net691;
 wire clknet_0_net619;
 wire clknet_1_0__leaf_net619;
 wire clknet_1_1__leaf_net619;
 wire clknet_0_net690;
 wire clknet_1_0__leaf_net690;
 wire clknet_1_1__leaf_net690;
 wire clknet_0_net689;
 wire clknet_1_0__leaf_net689;
 wire clknet_1_1__leaf_net689;
 wire clknet_0_net513;
 wire clknet_1_0__leaf_net513;
 wire clknet_1_1__leaf_net513;
 wire clknet_0_net672;
 wire clknet_1_0__leaf_net672;
 wire clknet_1_1__leaf_net672;
 wire clknet_0_net585;
 wire clknet_1_0__leaf_net585;
 wire clknet_1_1__leaf_net585;
 wire clknet_0_net597;
 wire clknet_1_0__leaf_net597;
 wire clknet_1_1__leaf_net597;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net586;
 wire clknet_1_0__leaf_net586;
 wire clknet_1_1__leaf_net586;
 wire clknet_0_net578;
 wire clknet_1_0__leaf_net578;
 wire clknet_1_1__leaf_net578;
 wire clknet_0_net476;
 wire clknet_1_0__leaf_net476;
 wire clknet_1_1__leaf_net476;
 wire clknet_0_net474;
 wire clknet_1_0__leaf_net474;
 wire clknet_1_1__leaf_net474;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net671;
 wire clknet_1_0__leaf_net671;
 wire clknet_1_1__leaf_net671;
 wire clknet_0_net670;
 wire clknet_1_0__leaf_net670;
 wire clknet_1_1__leaf_net670;
 wire clknet_0_net547;
 wire clknet_1_0__leaf_net547;
 wire clknet_1_1__leaf_net547;
 wire clknet_0_net794;
 wire clknet_1_0__leaf_net794;
 wire clknet_1_1__leaf_net794;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net530;
 wire clknet_1_0__leaf_net530;
 wire clknet_1_1__leaf_net530;
 wire clknet_0_net439;
 wire clknet_1_0__leaf_net439;
 wire clknet_1_1__leaf_net439;
 wire clknet_0_net643;
 wire clknet_1_0__leaf_net643;
 wire clknet_1_1__leaf_net643;
 wire clknet_0_net228;
 wire clknet_1_0__leaf_net228;
 wire clknet_1_1__leaf_net228;
 wire clknet_0_net238;
 wire clknet_1_0__leaf_net238;
 wire clknet_1_1__leaf_net238;
 wire clknet_0_net235;
 wire clknet_1_0__leaf_net235;
 wire clknet_1_1__leaf_net235;
 wire clknet_0_net241;
 wire clknet_1_0__leaf_net241;
 wire clknet_1_1__leaf_net241;
 wire clknet_0_net240;
 wire clknet_1_0__leaf_net240;
 wire clknet_1_1__leaf_net240;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net237;
 wire clknet_1_0__leaf_net237;
 wire clknet_1_1__leaf_net237;
 wire clknet_0_net249;
 wire clknet_1_0__leaf_net249;
 wire clknet_1_1__leaf_net249;
 wire clknet_0_net250;
 wire clknet_1_0__leaf_net250;
 wire clknet_1_1__leaf_net250;
 wire clknet_0_net236;
 wire clknet_1_0__leaf_net236;
 wire clknet_1_1__leaf_net236;
 wire clknet_0_net642;
 wire clknet_1_0__leaf_net642;
 wire clknet_1_1__leaf_net642;
 wire clknet_0_net143;
 wire clknet_1_0__leaf_net143;
 wire clknet_1_1__leaf_net143;
 wire clknet_0_net146;
 wire clknet_1_0__leaf_net146;
 wire clknet_1_1__leaf_net146;
 wire clknet_0_net815;
 wire clknet_1_0__leaf_net815;
 wire clknet_1_1__leaf_net815;
 wire clknet_0_net514;
 wire clknet_1_0__leaf_net514;
 wire clknet_1_1__leaf_net514;
 wire clknet_0_net835;
 wire clknet_1_0__leaf_net835;
 wire clknet_1_1__leaf_net835;
 wire clknet_0_net834;
 wire clknet_1_0__leaf_net834;
 wire clknet_1_1__leaf_net834;
 wire clknet_0_net145;
 wire clknet_1_0__leaf_net145;
 wire clknet_1_1__leaf_net145;
 wire clknet_0_net286;
 wire clknet_1_0__leaf_net286;
 wire clknet_1_1__leaf_net286;
 wire clknet_0_net165;
 wire clknet_1_0__leaf_net165;
 wire clknet_1_1__leaf_net165;
 wire clknet_0_net166;
 wire clknet_1_0__leaf_net166;
 wire clknet_1_1__leaf_net166;
 wire clknet_0_net796;
 wire clknet_1_0__leaf_net796;
 wire clknet_1_1__leaf_net796;
 wire clknet_0_net829;
 wire clknet_1_0__leaf_net829;
 wire clknet_1_1__leaf_net829;
 wire clknet_0_net852;
 wire clknet_1_0__leaf_net852;
 wire clknet_1_1__leaf_net852;
 wire clknet_0_net394;
 wire clknet_1_0__leaf_net394;
 wire clknet_1_1__leaf_net394;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire clknet_0_net169;
 wire clknet_1_0__leaf_net169;
 wire clknet_1_1__leaf_net169;
 wire clknet_0_net150;
 wire clknet_1_0__leaf_net150;
 wire clknet_1_1__leaf_net150;
 wire clknet_0_net843;
 wire clknet_1_0__leaf_net843;
 wire clknet_1_1__leaf_net843;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net378;
 wire clknet_1_0__leaf_net378;
 wire clknet_1_1__leaf_net378;
 wire clknet_0_net381;
 wire clknet_1_0__leaf_net381;
 wire clknet_1_1__leaf_net381;
 wire clknet_0_net379;
 wire clknet_1_0__leaf_net379;
 wire clknet_1_1__leaf_net379;
 wire clknet_0_net148;
 wire clknet_1_0__leaf_net148;
 wire clknet_1_1__leaf_net148;
 wire clknet_0_net155;
 wire clknet_1_0__leaf_net155;
 wire clknet_1_1__leaf_net155;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net164;
 wire clknet_1_0__leaf_net164;
 wire clknet_1_1__leaf_net164;
 wire clknet_0_net812;
 wire clknet_1_0__leaf_net812;
 wire clknet_1_1__leaf_net812;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net503;
 wire clknet_1_0__leaf_net503;
 wire clknet_1_1__leaf_net503;
 wire clknet_0_net501;
 wire clknet_1_0__leaf_net501;
 wire clknet_1_1__leaf_net501;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net491;
 wire clknet_1_0__leaf_net491;
 wire clknet_1_1__leaf_net491;
 wire clknet_0_net823;
 wire clknet_1_0__leaf_net823;
 wire clknet_1_1__leaf_net823;
 wire clknet_0_net261;
 wire clknet_1_0__leaf_net261;
 wire clknet_1_1__leaf_net261;
 wire clknet_0_net260;
 wire clknet_1_0__leaf_net260;
 wire clknet_1_1__leaf_net260;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net149;
 wire clknet_1_0__leaf_net149;
 wire clknet_1_1__leaf_net149;
 wire clknet_0_net147;
 wire clknet_1_0__leaf_net147;
 wire clknet_1_1__leaf_net147;
 wire clknet_0_net170;
 wire clknet_1_0__leaf_net170;
 wire clknet_1_1__leaf_net170;
 wire clknet_0_net848;
 wire clknet_1_0__leaf_net848;
 wire clknet_1_1__leaf_net848;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net818;
 wire clknet_1_0__leaf_net818;
 wire clknet_1_1__leaf_net818;
 wire clknet_0_net801;
 wire clknet_1_0__leaf_net801;
 wire clknet_1_1__leaf_net801;
 wire clknet_0_net144;
 wire clknet_1_0__leaf_net144;
 wire clknet_1_1__leaf_net144;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;

 sky130_fd_sc_hd__mux4_2 c100 (.A0(net23),
    .A1(net33),
    .A2(net34),
    .A3(net16),
    .S0(net35),
    .S1(net747),
    .X(net37));
 sky130_fd_sc_hd__nor2_4 c101 (.A(net739),
    .B(net33),
    .Y(net38));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net785),
    .A1(net37),
    .A2(net747),
    .A3(net38),
    .S0(net839),
    .S1(net13),
    .X(net39));
 sky130_fd_sc_hd__nor3b_4 c103 (.A(net37),
    .B(net39),
    .C_N(net839),
    .Y(net844));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net39),
    .A1(net35),
    .A2(net33),
    .A3(net844),
    .S0(net34),
    .S1(net38),
    .X(net40));
 sky130_fd_sc_hd__or2_1 c105 (.A(net12),
    .B(net844),
    .X(net41));
 sky130_fd_sc_hd__and2_1 c106 (.A(net771),
    .B(net839),
    .X(net42));
 sky130_fd_sc_hd__or2b_2 c107 (.A(net41),
    .B_N(net758),
    .X(net43));
 sky130_fd_sc_hd__or2_1 c108 (.A(net759),
    .B(net32),
    .X(net44));
 sky130_fd_sc_hd__nand2_1 c109 (.A(net11),
    .B(net844),
    .Y(net45));
 sky130_fd_sc_hd__and2b_1 c110 (.A_N(net43),
    .B(net844),
    .X(net46));
 sky130_fd_sc_hd__nand2_2 c111 (.A(net33),
    .B(net44),
    .Y(net47));
 sky130_fd_sc_hd__nand2b_1 c112 (.A_N(net760),
    .B(net33),
    .Y(net48));
 sky130_fd_sc_hd__and2_1 c113 (.A(net767),
    .B(net778),
    .X(net49));
 sky130_fd_sc_hd__nor2_1 c114 (.A(net758),
    .B(net47),
    .Y(net50));
 sky130_fd_sc_hd__nand2b_1 c115 (.A_N(net50),
    .B(net48),
    .Y(net51));
 sky130_fd_sc_hd__or4bb_2 c116 (.A(net51),
    .B(net8),
    .C_N(net49),
    .D_N(net32),
    .X(net52));
 sky130_fd_sc_hd__nand2b_1 c117 (.A_N(net49),
    .B(net52),
    .Y(net53));
 sky130_fd_sc_hd__and2_1 c118 (.A(net46),
    .B(net844),
    .X(net54));
 sky130_fd_sc_hd__or2_2 c119 (.A(net47),
    .B(net52),
    .X(net55));
 sky130_fd_sc_hd__mux4_4 c120 (.A0(net54),
    .A1(net55),
    .A2(net49),
    .A3(net50),
    .S0(net43),
    .S1(net44),
    .X(net56));
 sky130_fd_sc_hd__or2_1 c121 (.A(net48),
    .B(net49),
    .X(net57));
 sky130_fd_sc_hd__a2111o_2 c122 (.A1(net44),
    .A2(net47),
    .B1(net55),
    .C1(net43),
    .D1(net8),
    .X(net58));
 sky130_fd_sc_hd__or4bb_1 c123 (.A(net57),
    .B(net55),
    .C_N(net58),
    .D_N(net46),
    .X(net59));
 sky130_fd_sc_hd__mux4_4 c124 (.A0(net59),
    .A1(net52),
    .A2(net57),
    .A3(net54),
    .S0(net839),
    .S1(net897),
    .X(net60));
 sky130_fd_sc_hd__dfrbp_1 c125 (.CLK(clknet_leaf_13_clk),
    .D(net53),
    .RESET_B(net59),
    .Q(net62),
    .Q_N(net61));
 sky130_fd_sc_hd__nand2b_4 c126 (.A_N(net791),
    .B(net733),
    .Y(net63));
 sky130_fd_sc_hd__and3_1 c127 (.A(net742),
    .B(net755),
    .C(net735),
    .X(net64));
 sky130_fd_sc_hd__nor3b_1 c128 (.A(net745),
    .B(net788),
    .C_N(net735),
    .Y(net65));
 sky130_fd_sc_hd__mux4_2 c129 (.A0(net739),
    .A1(net733),
    .A2(net743),
    .A3(net735),
    .S0(net63),
    .S1(net895),
    .X(net66));
 sky130_fd_sc_hd__and3_2 c130 (.A(net65),
    .B(net740),
    .C(net895),
    .X(net67));
 sky130_fd_sc_hd__and3b_4 c131 (.A_N(net63),
    .B(net895),
    .C(net736),
    .X(net68));
 sky130_fd_sc_hd__and3_4 c132 (.A(net66),
    .B(net742),
    .C(net734),
    .X(net69));
 sky130_fd_sc_hd__nor3b_4 c133 (.A(net69),
    .B(net66),
    .C_N(net736),
    .Y(net70));
 sky130_fd_sc_hd__a2111oi_1 c134 (.A1(net63),
    .A2(net792),
    .B1(net737),
    .C1(net788),
    .D1(net895),
    .Y(net71));
 sky130_fd_sc_hd__nor3_2 c135 (.A(net791),
    .B(net961),
    .C(net64),
    .Y(net72));
 sky130_fd_sc_hd__o2111a_1 c136 (.A1(net792),
    .A2(net66),
    .B1(net72),
    .C1(net63),
    .D1(net68),
    .X(net73));
 sky130_fd_sc_hd__nand3_4 c137 (.A(net68),
    .B(net791),
    .C(net63),
    .Y(net74));
 sky130_fd_sc_hd__or2b_2 c138 (.A(net67),
    .B_N(net745),
    .X(net75));
 sky130_fd_sc_hd__or4bb_4 c139 (.A(net67),
    .B(net73),
    .C_N(net895),
    .D_N(net736),
    .X(net76));
 sky130_fd_sc_hd__nor3_4 c140 (.A(net735),
    .B(net742),
    .C(net70),
    .Y(net77));
 sky130_fd_sc_hd__nand3b_4 c141 (.A_N(net74),
    .B(net76),
    .C(net755),
    .Y(net78));
 sky130_fd_sc_hd__mux4_2 c142 (.A0(net69),
    .A1(net75),
    .A2(net78),
    .A3(net68),
    .S0(net66),
    .S1(net67),
    .X(net79));
 sky130_fd_sc_hd__nor3_1 c143 (.A(net79),
    .B(net67),
    .C(net77),
    .Y(net80));
 sky130_fd_sc_hd__a2111oi_2 c144 (.A1(net76),
    .A2(net78),
    .B1(net732),
    .C1(net75),
    .D1(net895),
    .Y(net81));
 sky130_fd_sc_hd__mux4_1 c145 (.A0(net80),
    .A1(net81),
    .A2(net75),
    .A3(net74),
    .S0(net66),
    .S1(net77),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c146 (.A0(net970),
    .A1(net82),
    .A2(net76),
    .A3(net894),
    .S0(net74),
    .S1(net895),
    .X(net83));
 sky130_fd_sc_hd__or4bb_2 c147 (.A(net757),
    .B(net740),
    .C_N(net759),
    .D_N(net900),
    .X(net84));
 sky130_fd_sc_hd__nand3b_2 c148 (.A_N(net64),
    .B(net736),
    .C(net83),
    .Y(net85));
 sky130_fd_sc_hd__or3b_1 c149 (.A(net882),
    .B(net788),
    .C_N(net895),
    .X(net86));
 sky130_fd_sc_hd__and3_1 c150 (.A(net70),
    .B(net750),
    .C(net902),
    .X(net87));
 sky130_fd_sc_hd__and2b_2 c151 (.A_N(net87),
    .B(net78),
    .X(net88));
 sky130_fd_sc_hd__or4bb_4 c152 (.A(net749),
    .B(net750),
    .C_N(net762),
    .D_N(net78),
    .X(net89));
 sky130_fd_sc_hd__and2_2 c153 (.A(net82),
    .B(net793),
    .X(net90));
 sky130_fd_sc_hd__mux4_2 c154 (.A0(net90),
    .A1(net884),
    .A2(net738),
    .A3(net86),
    .S0(net750),
    .S1(net768),
    .X(net91));
 sky130_fd_sc_hd__nor2_1 c155 (.A(net761),
    .B(net90),
    .Y(net92));
 sky130_fd_sc_hd__or2_1 c156 (.A(net83),
    .B(net90),
    .X(net93));
 sky130_fd_sc_hd__nand3b_1 c157 (.A_N(net93),
    .B(net882),
    .C(net85),
    .Y(net94));
 sky130_fd_sc_hd__nand3b_1 c158 (.A_N(net753),
    .B(net92),
    .C(net91),
    .Y(net95));
 sky130_fd_sc_hd__a2111oi_4 c159 (.A1(net736),
    .A2(net89),
    .B1(net90),
    .C1(net94),
    .D1(net880),
    .Y(net96));
 sky130_fd_sc_hd__nor2_4 c160 (.A(net737),
    .B(net92),
    .Y(net97));
 sky130_fd_sc_hd__o2111a_2 c161 (.A1(net95),
    .A2(net97),
    .B1(net78),
    .C1(net753),
    .D1(net81),
    .X(net98));
 sky130_fd_sc_hd__and3_1 c162 (.A(net98),
    .B(net736),
    .C(net95),
    .X(net99));
 sky130_fd_sc_hd__or4bb_4 c163 (.A(net99),
    .B(net98),
    .C_N(net895),
    .D_N(net88),
    .X(net100));
 sky130_fd_sc_hd__sdfrbp_1 c164 (.CLK(clknet_leaf_6_clk),
    .D(net96),
    .RESET_B(net754),
    .SCD(net100),
    .SCE(net90),
    .Q(net102),
    .Q_N(net101));
 sky130_fd_sc_hd__mux4_1 c165 (.A0(net92),
    .A1(net100),
    .A2(net98),
    .A3(net97),
    .S0(net91),
    .S1(net70),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net94),
    .A1(net89),
    .A2(net91),
    .A3(net90),
    .S0(net98),
    .S1(net915),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 c167 (.A0(net94),
    .A1(net100),
    .A2(net95),
    .A3(net96),
    .S0(net74),
    .S1(net915),
    .X(net105));
 sky130_fd_sc_hd__nand3_1 c168 (.A(net75),
    .B(net770),
    .C(net101),
    .Y(net106));
 sky130_fd_sc_hd__nor2b_1 c169 (.A(net79),
    .B_N(net788),
    .Y(net107));
 sky130_fd_sc_hd__or3_1 c170 (.A(net104),
    .B(net106),
    .C(net78),
    .X(net108));
 sky130_fd_sc_hd__sdfrbp_1 c171 (.CLK(clknet_leaf_6_clk),
    .D(net770),
    .RESET_B(net108),
    .SCD(net75),
    .SCE(net779),
    .Q(net110),
    .Q_N(net109));
 sky130_fd_sc_hd__nor3b_1 c172 (.A(net102),
    .B(net107),
    .C_N(net784),
    .Y(net111));
 sky130_fd_sc_hd__and2b_1 c173 (.A_N(net106),
    .B(net107),
    .X(net112));
 sky130_fd_sc_hd__and2_1 c174 (.A(net78),
    .B(net111),
    .X(net113));
 sky130_fd_sc_hd__and2_2 c175 (.A(net111),
    .B(net783),
    .X(net114));
 sky130_fd_sc_hd__nand2b_1 c176 (.A_N(net894),
    .B(net113),
    .Y(net115));
 sky130_fd_sc_hd__mux4_1 c177 (.A0(net110),
    .A1(net106),
    .A2(net75),
    .A3(net878),
    .S0(net79),
    .S1(net882),
    .X(net116));
 sky130_fd_sc_hd__dfbbn_1 c178 (.CLK_N(clknet_leaf_6_clk),
    .D(net108),
    .RESET_B(net878),
    .SET_B(net114),
    .Q(net118),
    .Q_N(net117));
 sky130_fd_sc_hd__nand3b_4 c179 (.A_N(net733),
    .B(net752),
    .C(net102),
    .Y(net119));
 sky130_fd_sc_hd__mux4_2 c180 (.A0(net116),
    .A1(net96),
    .A2(net91),
    .A3(net117),
    .S0(net109),
    .S1(net114),
    .X(net120));
 sky130_fd_sc_hd__or3b_4 c181 (.A(net120),
    .B(net106),
    .C_N(net115),
    .X(net121));
 sky130_fd_sc_hd__sdfbbn_1 c182 (.CLK_N(clknet_leaf_6_clk),
    .D(net113),
    .RESET_B(net121),
    .SCD(net120),
    .SCE(net112),
    .SET_B(net779),
    .Q(net123),
    .Q_N(net122));
 sky130_fd_sc_hd__sdfbbn_1 c183 (.CLK_N(clknet_leaf_7_clk),
    .D(net923),
    .RESET_B(net120),
    .SCD(net114),
    .SCE(net116),
    .SET_B(net121),
    .Q(net125),
    .Q_N(net124));
 sky130_fd_sc_hd__mux4_4 c184 (.A0(net115),
    .A1(net120),
    .A2(net111),
    .A3(net96),
    .S0(net783),
    .S1(net121),
    .X(net126));
 sky130_fd_sc_hd__dfbbn_2 c185 (.CLK_N(clknet_leaf_7_clk),
    .D(net121),
    .RESET_B(net940),
    .SET_B(net641),
    .Q(net128),
    .Q_N(net127));
 sky130_fd_sc_hd__mux4_1 c186 (.A0(net769),
    .A1(net121),
    .A2(net112),
    .A3(net127),
    .S0(net124),
    .S1(net641),
    .X(net129));
 sky130_fd_sc_hd__mux4_4 c187 (.A0(net107),
    .A1(net114),
    .A2(net783),
    .A3(net0),
    .S0(net641),
    .S1(clknet_1_0__leaf_net642),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net130),
    .A1(net108),
    .A2(net128),
    .A3(net122),
    .S0(net120),
    .S1(net641),
    .X(net131));
 sky130_fd_sc_hd__nor2b_1 c189 (.A(net10),
    .B_N(net19),
    .Y(net132));
 sky130_fd_sc_hd__sdfrtn_1 c190 (.CLK_N(clknet_leaf_7_clk),
    .D(net750),
    .RESET_B(net10),
    .SCD(net121),
    .SCE(clknet_1_1__leaf_net642),
    .Q(net133));
 sky130_fd_sc_hd__a2111oi_1 c191 (.A1(net773),
    .A2(net0),
    .B1(net133),
    .C1(net897),
    .D1(net732),
    .Y(net134));
 sky130_fd_sc_hd__nand2b_4 c192 (.A_N(net15),
    .B(net20),
    .Y(net135));
 sky130_fd_sc_hd__nand3b_1 c193 (.A_N(net19),
    .B(net125),
    .C(net135),
    .Y(net136));
 sky130_fd_sc_hd__nor2b_2 c194 (.A(net887),
    .B_N(net88),
    .Y(net137));
 sky130_fd_sc_hd__o2111ai_4 c195 (.A1(net0),
    .A2(net21),
    .B1(net137),
    .C1(net74),
    .D1(net135),
    .Y(net138));
 sky130_fd_sc_hd__and3b_4 c196 (.A_N(net755),
    .B(net19),
    .C(net10),
    .X(net139));
 sky130_fd_sc_hd__nor3_1 c197 (.A(net783),
    .B(net134),
    .C(net899),
    .Y(net140));
 sky130_fd_sc_hd__a2111o_1 c198 (.A1(net133),
    .A2(net74),
    .B1(net773),
    .C1(net135),
    .D1(net139),
    .X(net141));
 sky130_fd_sc_hd__or4bb_4 c199 (.A(net88),
    .B(net135),
    .C_N(clknet_1_0__leaf_net642),
    .D_N(net139),
    .X(net142));
 sky130_fd_sc_hd__or4bb_4 c200 (.A(net135),
    .B(net968),
    .C_N(clknet_1_1__leaf_net642),
    .D_N(clknet_1_1__leaf_net142),
    .X(net143));
 sky130_fd_sc_hd__o2111a_2 c201 (.A1(net139),
    .A2(net135),
    .B1(net15),
    .C1(net141),
    .D1(clknet_1_1__leaf_net142),
    .X(net144));
 sky130_fd_sc_hd__mux4_2 c202 (.A0(net132),
    .A1(net21),
    .A2(net135),
    .A3(net138),
    .S0(clknet_1_1__leaf_net143),
    .S1(clknet_1_1__leaf_net142),
    .X(net145));
 sky130_fd_sc_hd__or4bb_2 c203 (.A(clknet_1_0__leaf_net143),
    .B(net899),
    .C_N(net124),
    .D_N(net976),
    .X(net146));
 sky130_fd_sc_hd__nand3_4 c204 (.A(net136),
    .B(net15),
    .C(clknet_1_1__leaf_net142),
    .Y(net147));
 sky130_fd_sc_hd__mux4_2 c205 (.A0(net138),
    .A1(net135),
    .A2(clknet_1_1__leaf_net144),
    .A3(clknet_1_0__leaf_net145),
    .S0(net14),
    .S1(net127),
    .X(net148));
 sky130_fd_sc_hd__mux4_4 c206 (.A0(net141),
    .A1(net140),
    .A2(net125),
    .A3(clknet_1_1__leaf_net146),
    .S0(net899),
    .S1(net905),
    .X(net834));
 sky130_fd_sc_hd__and3_2 c207 (.A(net21),
    .B(net139),
    .C(clknet_1_1__leaf_net142),
    .X(net149));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(clknet_1_0__leaf_net144),
    .A1(clknet_1_1__leaf_net149),
    .A2(net132),
    .A3(net135),
    .S0(net899),
    .S1(net977),
    .X(net843));
 sky130_fd_sc_hd__mux4_4 c209 (.A0(clknet_1_0__leaf_net149),
    .A1(net977),
    .A2(net138),
    .A3(net135),
    .S0(net976),
    .S1(net899),
    .X(net150));
 sky130_fd_sc_hd__mux4_2 c210 (.A0(net31),
    .A1(net34),
    .A2(net14),
    .A3(clknet_1_0__leaf_net148),
    .S0(clknet_1_1__leaf_net146),
    .S1(net25),
    .X(net815));
 sky130_fd_sc_hd__nand2b_1 c211 (.A_N(net26),
    .B(net8),
    .Y(net151));
 sky130_fd_sc_hd__or2b_2 c212 (.A(net140),
    .B_N(net137),
    .X(net152));
 sky130_fd_sc_hd__nor2b_1 c213 (.A(net152),
    .B_N(net74),
    .Y(net153));
 sky130_fd_sc_hd__nand2b_1 c214 (.A_N(net137),
    .B(net97),
    .Y(net154));
 sky130_fd_sc_hd__nand3b_4 c215 (.A_N(clknet_1_1__leaf_net148),
    .B(net97),
    .C(net38),
    .Y(net155));
 sky130_fd_sc_hd__a2111oi_4 c216 (.A1(net879),
    .A2(net766),
    .B1(net38),
    .C1(net844),
    .D1(clknet_1_1__leaf_net145),
    .Y(net156));
 sky130_fd_sc_hd__a2111o_1 c217 (.A1(net88),
    .A2(net128),
    .B1(net137),
    .C1(net8),
    .D1(net152),
    .X(net157));
 sky130_fd_sc_hd__and3b_1 c218 (.A_N(net25),
    .B(net137),
    .C(net777),
    .X(net158));
 sky130_fd_sc_hd__and3_1 c219 (.A(net151),
    .B(net25),
    .C(net782),
    .X(net159));
 sky130_fd_sc_hd__nor3b_1 c220 (.A(net35),
    .B(clknet_1_0__leaf_net147),
    .C_N(net27),
    .Y(net160));
 sky130_fd_sc_hd__nor2b_1 c221 (.A(net158),
    .B_N(net27),
    .Y(net161));
 sky130_fd_sc_hd__or2_1 c222 (.A(clknet_1_0__leaf_net160),
    .B(net152),
    .X(net818));
 sky130_fd_sc_hd__nor3_4 c223 (.A(net97),
    .B(net766),
    .C(net784),
    .Y(net849));
 sky130_fd_sc_hd__and2b_2 c224 (.A_N(net125),
    .B(clknet_1_1__leaf_net155),
    .X(net162));
 sky130_fd_sc_hd__mux4_2 c225 (.A0(net766),
    .A1(net161),
    .A2(net735),
    .A3(net38),
    .S0(net849),
    .S1(net36),
    .X(net163));
 sky130_fd_sc_hd__o2111ai_4 c226 (.A1(clknet_1_1__leaf_net162),
    .A2(net972),
    .B1(clknet_1_0__leaf_net147),
    .C1(net40),
    .D1(net31),
    .Y(net812));
 sky130_fd_sc_hd__nand3b_1 c227 (.A_N(net74),
    .B(clknet_1_0__leaf_net162),
    .C(clknet_1_0__leaf_net160),
    .Y(net164));
 sky130_fd_sc_hd__and2b_1 c228 (.A_N(net153),
    .B(clknet_1_0__leaf_net145),
    .X(net165));
 sky130_fd_sc_hd__and3b_2 c229 (.A_N(clknet_1_0__leaf_net165),
    .B(clknet_1_1__leaf_net160),
    .C(clknet_1_0__leaf_net818),
    .X(net829));
 sky130_fd_sc_hd__mux4_4 c230 (.A0(net30),
    .A1(net138),
    .A2(net97),
    .A3(clknet_1_1__leaf_net165),
    .S0(clknet_1_1__leaf_net829),
    .S1(net25),
    .X(net166));
 sky130_fd_sc_hd__nor3b_2 c231 (.A(net52),
    .B(net849),
    .C_N(net43),
    .Y(net825));
 sky130_fd_sc_hd__or3b_1 c232 (.A(net42),
    .B(clknet_1_0__leaf_net156),
    .C_N(net849),
    .X(net167));
 sky130_fd_sc_hd__nand3b_2 c233 (.A_N(clknet_1_1__leaf_net147),
    .B(net138),
    .C(net638),
    .Y(net848));
 sky130_fd_sc_hd__nand3_2 c234 (.A(clknet_1_0__leaf_net166),
    .B(clknet_1_1__leaf_net834),
    .C(net847),
    .Y(net168));
 sky130_fd_sc_hd__o2111a_1 c235 (.A1(clknet_1_1__leaf_net156),
    .A2(net825),
    .B1(net58),
    .C1(net47),
    .D1(net8),
    .X(net169));
 sky130_fd_sc_hd__or4bb_1 c236 (.A(net43),
    .B(clknet_1_0__leaf_net147),
    .C_N(net161),
    .D_N(net32),
    .X(net170));
 sky130_fd_sc_hd__a2111oi_1 c237 (.A1(net62),
    .A2(net49),
    .B1(net58),
    .C1(net42),
    .D1(net638),
    .Y(net171));
 sky130_fd_sc_hd__and3b_4 c238 (.A_N(clknet_1_1__leaf_net170),
    .B(clknet_1_0__leaf_net848),
    .C(net52),
    .X(net172));
 sky130_fd_sc_hd__nor3_1 c239 (.A(net32),
    .B(clknet_1_1__leaf_net166),
    .C(clknet_1_0__leaf_net170),
    .Y(net796));
 sky130_fd_sc_hd__sdfbbp_1 c240 (.CLK(clknet_leaf_15_clk),
    .D(net902),
    .RESET_B(net759),
    .SCD(clknet_1_0__leaf_net796),
    .SCE(clknet_1_0__leaf_net812),
    .SET_B(net161),
    .Q(net174),
    .Q_N(net173));
 sky130_fd_sc_hd__sdfbbn_1 c241 (.CLK_N(clknet_leaf_14_clk),
    .D(net161),
    .RESET_B(clknet_1_1__leaf_net812),
    .SCD(clknet_1_1__leaf_net818),
    .SCE(net844),
    .SET_B(net173),
    .Q(net810),
    .Q_N(net175));
 sky130_fd_sc_hd__sdfrtp_1 c242 (.CLK(clknet_leaf_15_clk),
    .D(net174),
    .RESET_B(net825),
    .SCD(clknet_1_1__leaf_net796),
    .SCE(net175),
    .Q(net831));
 sky130_fd_sc_hd__o2111ai_4 c243 (.A1(net55),
    .A2(net47),
    .B1(net934),
    .C1(net782),
    .D1(net138),
    .Y(net176));
 sky130_fd_sc_hd__mux4_4 c244 (.A0(net172),
    .A1(clknet_1_0__leaf_net169),
    .A2(clknet_1_1__leaf_net843),
    .A3(clknet_1_1__leaf_net147),
    .S0(net42),
    .S1(clknet_1_1__leaf_net818),
    .X(net177));
 sky130_fd_sc_hd__a2111o_4 c245 (.A1(net735),
    .A2(net810),
    .B1(net902),
    .C1(clknet_1_1__leaf_net147),
    .D1(net824),
    .X(net842));
 sky130_fd_sc_hd__dfbbp_1 c246 (.CLK(clknet_leaf_13_clk),
    .D(net168),
    .RESET_B(clknet_1_0__leaf_net848),
    .SET_B(net637),
    .Q(net821),
    .Q_N(net178));
 sky130_fd_sc_hd__sdfbbn_1 c247 (.CLK_N(clknet_leaf_14_clk),
    .D(net45),
    .RESET_B(net821),
    .SCD(net175),
    .SCE(net61),
    .SET_B(clknet_1_1__leaf_net169),
    .Q(net845),
    .Q_N(net179));
 sky130_fd_sc_hd__or4bb_1 c248 (.A(net167),
    .B(net845),
    .C_N(net55),
    .D_N(net45),
    .X(net180));
 sky130_fd_sc_hd__sdfbbp_1 c249 (.CLK(clknet_leaf_13_clk),
    .D(net171),
    .RESET_B(net43),
    .SCD(net845),
    .SCE(net935),
    .SET_B(net176),
    .Q(net820));
 sky130_fd_sc_hd__sdfrtp_1 c250 (.CLK(clknet_leaf_14_clk),
    .D(net180),
    .RESET_B(clknet_1_0__leaf_net796),
    .SCD(net174),
    .SCE(net179),
    .Q(net181));
 sky130_fd_sc_hd__and3_1 c251 (.A(net181),
    .B(net902),
    .C(net179),
    .X(net182));
 sky130_fd_sc_hd__nor2b_1 c252 (.A(net735),
    .B_N(net68),
    .Y(net183));
 sky130_fd_sc_hd__or4bb_4 c253 (.A(net77),
    .B(net792),
    .C_N(net788),
    .D_N(net69),
    .X(net184));
 sky130_fd_sc_hd__and2b_1 c254 (.A_N(net183),
    .B(net77),
    .X(net185));
 sky130_fd_sc_hd__or2_4 c255 (.A(net67),
    .B(net744),
    .X(net186));
 sky130_fd_sc_hd__nor2b_2 c256 (.A(net185),
    .B_N(net186),
    .Y(net187));
 sky130_fd_sc_hd__nor2b_2 c257 (.A(net777),
    .B_N(net183),
    .Y(net188));
 sky130_fd_sc_hd__or2_1 c258 (.A(net187),
    .B(net883),
    .X(net189));
 sky130_fd_sc_hd__o2111ai_4 c259 (.A1(net77),
    .A2(net69),
    .B1(net890),
    .C1(net184),
    .D1(net68),
    .Y(net190));
 sky130_fd_sc_hd__or4bb_4 c260 (.A(net743),
    .B(net184),
    .C_N(net67),
    .D_N(net896),
    .X(net827));
 sky130_fd_sc_hd__mux4_2 c261 (.A0(net73),
    .A1(net189),
    .A2(net187),
    .A3(net184),
    .S0(net186),
    .S1(net883),
    .X(net191));
 sky130_fd_sc_hd__nor3_1 c262 (.A(net183),
    .B(net190),
    .C(net186),
    .Y(net192));
 sky130_fd_sc_hd__a2111oi_1 c263 (.A1(net186),
    .A2(net744),
    .B1(net184),
    .C1(net877),
    .D1(net732),
    .Y(net193));
 sky130_fd_sc_hd__o2111a_1 c264 (.A1(net189),
    .A2(net184),
    .B1(net876),
    .C1(net877),
    .D1(net190),
    .X(net194));
 sky130_fd_sc_hd__mux4_2 c265 (.A0(net745),
    .A1(net735),
    .A2(net77),
    .A3(net788),
    .S0(net184),
    .S1(net187),
    .X(net195));
 sky130_fd_sc_hd__or2_2 c266 (.A(net734),
    .B(net194),
    .X(net196));
 sky130_fd_sc_hd__mux4_2 c267 (.A0(net195),
    .A1(net194),
    .A2(net877),
    .A3(net743),
    .S0(net189),
    .S1(net183),
    .X(net197));
 sky130_fd_sc_hd__or3_4 c268 (.A(net827),
    .B(net876),
    .C(net883),
    .X(net198));
 sky130_fd_sc_hd__mux4_2 c269 (.A0(net192),
    .A1(net187),
    .A2(net67),
    .A3(net827),
    .S0(net195),
    .S1(net196),
    .X(net199));
 sky130_fd_sc_hd__and2_2 c270 (.A(net197),
    .B(net72),
    .X(net795));
 sky130_fd_sc_hd__mux4_1 c271 (.A0(net193),
    .A1(net199),
    .A2(net883),
    .A3(net196),
    .S0(net187),
    .S1(net877),
    .X(net200));
 sky130_fd_sc_hd__nor3b_1 c272 (.A(net199),
    .B(net186),
    .C_N(net197),
    .Y(net201));
 sky130_fd_sc_hd__nor2b_1 c273 (.A(net901),
    .B_N(net827),
    .Y(net202));
 sky130_fd_sc_hd__nor2b_1 c274 (.A(net884),
    .B_N(net866),
    .Y(net203));
 sky130_fd_sc_hd__and2_1 c275 (.A(net744),
    .B(net793),
    .X(net204));
 sky130_fd_sc_hd__dfrbp_2 c276 (.CLK(clknet_leaf_8_clk),
    .D(net754),
    .RESET_B(net100),
    .Q(net206),
    .Q_N(net205));
 sky130_fd_sc_hd__nand2b_1 c277 (.A_N(net89),
    .B(net738),
    .Y(net207));
 sky130_fd_sc_hd__and2_1 c278 (.A(net204),
    .B(net76),
    .X(net208));
 sky130_fd_sc_hd__or2_4 c279 (.A(net207),
    .B(net89),
    .X(net209));
 sky130_fd_sc_hd__nand2b_1 c280 (.A_N(net793),
    .B(net204),
    .Y(net210));
 sky130_fd_sc_hd__or4bb_1 c281 (.A(net210),
    .B(net900),
    .C_N(net190),
    .D_N(net895),
    .X(net211));
 sky130_fd_sc_hd__a2111o_4 c282 (.A1(net190),
    .A2(net209),
    .B1(net208),
    .C1(net748),
    .D1(net640),
    .X(net212));
 sky130_fd_sc_hd__or4bb_1 c283 (.A(net208),
    .B(net900),
    .C_N(net206),
    .D_N(net211),
    .X(net213));
 sky130_fd_sc_hd__or3_1 c284 (.A(net208),
    .B(net188),
    .C(net205),
    .X(net214));
 sky130_fd_sc_hd__sdfrtp_4 c285 (.CLK(clknet_leaf_5_clk),
    .D(net211),
    .RESET_B(net202),
    .SCD(net100),
    .SCE(net795),
    .Q(net215));
 sky130_fd_sc_hd__mux4_4 c286 (.A0(net215),
    .A1(net204),
    .A2(net212),
    .A3(net209),
    .S0(net100),
    .S1(net210),
    .X(net216));
 sky130_fd_sc_hd__and2b_1 c287 (.A_N(net203),
    .B(net89),
    .X(net217));
 sky130_fd_sc_hd__sdfbbn_1 c288 (.CLK_N(clknet_leaf_5_clk),
    .D(net100),
    .RESET_B(net203),
    .SCD(net212),
    .SCE(net89),
    .SET_B(net198),
    .Q(net219),
    .Q_N(net218));
 sky130_fd_sc_hd__nor2_4 c289 (.A(net219),
    .B(net209),
    .Y(net220));
 sky130_fd_sc_hd__mux4_2 c290 (.A0(net214),
    .A1(net209),
    .A2(net884),
    .A3(net202),
    .S0(net212),
    .S1(net644),
    .X(net221));
 sky130_fd_sc_hd__a2111oi_1 c291 (.A1(net214),
    .A2(net219),
    .B1(net207),
    .C1(net884),
    .D1(net877),
    .Y(net222));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net222),
    .A1(net215),
    .A2(net884),
    .A3(net196),
    .S0(net217),
    .S1(net645),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net217),
    .A1(net214),
    .A2(net218),
    .A3(net957),
    .S0(net215),
    .S1(net809),
    .X(net224));
 sky130_fd_sc_hd__nand3b_4 c294 (.A_N(net788),
    .B(net119),
    .C(clknet_1_0__leaf_net643),
    .Y(net225));
 sky130_fd_sc_hd__nand3b_4 c295 (.A_N(net786),
    .B(net122),
    .C(net205),
    .Y(net226));
 sky130_fd_sc_hd__nor2_1 c296 (.A(net196),
    .B(net647),
    .Y(net227));
 sky130_fd_sc_hd__and2_0 c297 (.A(net119),
    .B(clknet_1_1__leaf_net643),
    .X(net228));
 sky130_fd_sc_hd__mux4_2 c298 (.A0(net114),
    .A1(net227),
    .A2(clknet_1_0__leaf_net228),
    .A3(net226),
    .S0(net752),
    .S1(net896),
    .X(net229));
 sky130_fd_sc_hd__or4bb_1 c299 (.A(net779),
    .B(net206),
    .C_N(net123),
    .D_N(net648),
    .X(net230));
 sky130_fd_sc_hd__or2_1 c300 (.A(net787),
    .B(net746),
    .X(net231));
 sky130_fd_sc_hd__nor2b_1 c301 (.A(net91),
    .B_N(net227),
    .Y(net232));
 sky130_fd_sc_hd__and3b_2 c302 (.A_N(net231),
    .B(net98),
    .C(net226),
    .X(net233));
 sky130_fd_sc_hd__nand2_4 c303 (.A(net226),
    .B(net114),
    .Y(net234));
 sky130_fd_sc_hd__nand3b_4 c304 (.A_N(net225),
    .B(net234),
    .C(net215),
    .Y(net235));
 sky130_fd_sc_hd__or3_4 c305 (.A(clknet_1_0__leaf_net235),
    .B(net212),
    .C(net779),
    .X(net236));
 sky130_fd_sc_hd__nand3b_1 c306 (.A_N(net756),
    .B(net234),
    .C(clknet_1_0__leaf_net235),
    .Y(net237));
 sky130_fd_sc_hd__nor3b_1 c307 (.A(net229),
    .B(clknet_1_0__leaf_net235),
    .C_N(net875),
    .Y(net238));
 sky130_fd_sc_hd__nor2_1 c308 (.A(net230),
    .B(net127),
    .Y(net239));
 sky130_fd_sc_hd__and2_2 c309 (.A(clknet_1_1__leaf_net236),
    .B(clknet_1_1__leaf_net235),
    .X(net240));
 sky130_fd_sc_hd__nand3_4 c310 (.A(net226),
    .B(clknet_1_1__leaf_net235),
    .C(net233),
    .Y(net241));
 sky130_fd_sc_hd__mux4_4 c311 (.A0(net233),
    .A1(clknet_1_1__leaf_net241),
    .A2(net119),
    .A3(clknet_1_1__leaf_net240),
    .S0(net98),
    .S1(clknet_1_0__leaf_net236),
    .X(net242));
 sky130_fd_sc_hd__mux4_2 c312 (.A0(net239),
    .A1(clknet_1_1__leaf_net235),
    .A2(clknet_1_0__leaf_net241),
    .A3(net234),
    .S0(net827),
    .S1(net892),
    .X(net243));
 sky130_fd_sc_hd__sdfsbp_1 c313 (.CLK(clknet_leaf_8_clk),
    .D(net232),
    .SCD(clknet_1_1__leaf_net241),
    .SCE(net892),
    .SET_B(net649),
    .Q(net245),
    .Q_N(net244));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net232),
    .A1(clknet_1_1__leaf_net240),
    .A2(clknet_1_0__leaf_net237),
    .A3(net233),
    .S0(net892),
    .S1(net649),
    .X(net246));
 sky130_fd_sc_hd__sdfsbp_1 c315 (.CLK(clknet_leaf_9_clk),
    .D(net231),
    .SCD(clknet_1_0__leaf_net146),
    .SCE(net121),
    .SET_B(net905),
    .Q(net248),
    .Q_N(net247));
 sky130_fd_sc_hd__or4bb_4 c316 (.A(clknet_1_1__leaf_net237),
    .B(net20),
    .C_N(net245),
    .D_N(net905),
    .X(net249));
 sky130_fd_sc_hd__a2111oi_4 c317 (.A1(clknet_1_1__leaf_net249),
    .A2(net119),
    .B1(net827),
    .C1(net244),
    .D1(net646),
    .Y(net250));
 sky130_fd_sc_hd__sdfxbp_1 c318 (.CLK(clknet_leaf_11_clk),
    .D(clknet_1_1__leaf_net150),
    .SCD(clknet_1_1__leaf_net228),
    .SCE(clknet_1_1__leaf_net250),
    .Q(net252),
    .Q_N(net251));
 sky130_fd_sc_hd__sdfxbp_1 c319 (.CLK(clknet_leaf_11_clk),
    .D(clknet_1_0__leaf_net250),
    .SCD(clknet_1_0__leaf_net834),
    .SCE(net932),
    .Q(net254),
    .Q_N(net253));
 sky130_fd_sc_hd__nor3_1 c320 (.A(net245),
    .B(net248),
    .C(clknet_1_0__leaf_net843),
    .Y(net255));
 sky130_fd_sc_hd__and3b_4 c321 (.A_N(net20),
    .B(net882),
    .C(net244),
    .X(net256));
 sky130_fd_sc_hd__sdfxtp_1 c322 (.CLK(clknet_leaf_8_clk),
    .D(clknet_1_0__leaf_net241),
    .SCD(net938),
    .SCE(net221),
    .Q(net257));
 sky130_fd_sc_hd__nor3_1 c323 (.A(clknet_1_1__leaf_net255),
    .B(clknet_1_0__leaf_net249),
    .C(clknet_1_0__leaf_net843),
    .Y(net258));
 sky130_fd_sc_hd__sdfxtp_1 c324 (.CLK(clknet_leaf_8_clk),
    .D(net928),
    .SCD(clknet_1_0__leaf_net146),
    .SCE(clknet_1_0__leaf_net241),
    .Q(net259));
 sky130_fd_sc_hd__or4bb_2 c325 (.A(net932),
    .B(net865),
    .C_N(net875),
    .D_N(net976),
    .X(net260));
 sky130_fd_sc_hd__a2111oi_1 c326 (.A1(net259),
    .A2(clknet_1_1__leaf_net260),
    .B1(net253),
    .C1(net898),
    .D1(net905),
    .Y(net261));
 sky130_fd_sc_hd__sdfbbn_1 c327 (.CLK_N(clknet_leaf_10_clk),
    .D(net875),
    .RESET_B(net827),
    .SCD(net259),
    .SCE(clknet_1_1__leaf_net261),
    .SET_B(net257),
    .Q(net830),
    .Q_N(net262));
 sky130_fd_sc_hd__mux4_2 c328 (.A0(net258),
    .A1(clknet_1_0__leaf_net228),
    .A2(net257),
    .A3(clknet_1_0__leaf_net260),
    .S0(net978),
    .S1(net220),
    .X(net263));
 sky130_fd_sc_hd__sdfbbp_1 c329 (.CLK(clknet_leaf_10_clk),
    .D(clknet_1_0__leaf_net260),
    .RESET_B(net875),
    .SCD(net18),
    .SCE(clknet_1_1__leaf_net261),
    .SET_B(clknet_1_0__leaf_net843),
    .Q(net265),
    .Q_N(net264));
 sky130_fd_sc_hd__mux4_2 c330 (.A0(net256),
    .A1(clknet_1_0__leaf_net150),
    .A2(net233),
    .A3(clknet_1_0__leaf_net145),
    .S0(net648),
    .S1(net650),
    .X(net266));
 sky130_fd_sc_hd__sdfbbn_1 c331 (.CLK_N(clknet_leaf_10_clk),
    .D(net266),
    .RESET_B(net8),
    .SCD(net256),
    .SCE(net264),
    .SET_B(clknet_1_1__leaf_net261),
    .Q(net268),
    .Q_N(net267));
 sky130_fd_sc_hd__nand3_4 c332 (.A(net267),
    .B(clknet_1_1__leaf_net260),
    .C(net650),
    .Y(net269));
 sky130_fd_sc_hd__sdfbbn_1 c333 (.CLK_N(clknet_leaf_10_clk),
    .D(net925),
    .RESET_B(clknet_1_1__leaf_net261),
    .SCD(net254),
    .SCE(net245),
    .SET_B(clknet_1_0__leaf_net146),
    .Q(net271),
    .Q_N(net270));
 sky130_fd_sc_hd__mux4_4 c334 (.A0(clknet_1_0__leaf_net250),
    .A1(net265),
    .A2(net259),
    .A3(clknet_1_0__leaf_net261),
    .S0(net270),
    .S1(clknet_1_0__leaf_net269),
    .X(net272));
 sky130_fd_sc_hd__mux4_2 c335 (.A0(net254),
    .A1(net271),
    .A2(clknet_1_0__leaf_net269),
    .A3(net264),
    .S0(net782),
    .S1(net891),
    .X(net273));
 sky130_fd_sc_hd__and3_1 c336 (.A(net40),
    .B(net271),
    .C(net891),
    .X(net274));
 sky130_fd_sc_hd__sdfxtp_1 c337 (.CLK(clknet_leaf_11_clk),
    .D(net157),
    .SCD(clknet_1_0__leaf_net164),
    .SCE(clknet_1_1__leaf_net236),
    .Q(net275));
 sky130_fd_sc_hd__nor3b_1 c338 (.A(net38),
    .B(net839),
    .C_N(net40),
    .Y(net276));
 sky130_fd_sc_hd__nand3_4 c339 (.A(net128),
    .B(net275),
    .C(net205),
    .Y(net832));
 sky130_fd_sc_hd__or3b_1 c340 (.A(net14),
    .B(net274),
    .C_N(net782),
    .X(net277));
 sky130_fd_sc_hd__nand3_1 c341 (.A(clknet_1_1__leaf_net146),
    .B(net38),
    .C(net251),
    .Y(net278));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net154),
    .A1(net277),
    .A2(net275),
    .A3(net262),
    .S0(net832),
    .S1(net651),
    .X(net279));
 sky130_fd_sc_hd__nor3_1 c343 (.A(net277),
    .B(net233),
    .C(net275),
    .Y(net850));
 sky130_fd_sc_hd__dfbbn_1 c344 (.CLK_N(clknet_leaf_11_clk),
    .D(clknet_1_1__leaf_net164),
    .RESET_B(net262),
    .SET_B(clknet_1_0__leaf_net815),
    .Q(net281),
    .Q_N(net280));
 sky130_fd_sc_hd__sdfstp_1 c345 (.CLK(clknet_leaf_18_clk),
    .D(net121),
    .SCD(net276),
    .SCE(net827),
    .SET_B(net892),
    .Q(net282));
 sky130_fd_sc_hd__nand2b_1 c346 (.A_N(net274),
    .B(net206),
    .Y(net840));
 sky130_fd_sc_hd__dfbbn_1 c347 (.CLK_N(clknet_leaf_15_clk),
    .D(net921),
    .RESET_B(net275),
    .SET_B(clknet_1_1__leaf_net238),
    .Q(net283));
 sky130_fd_sc_hd__sdfstp_1 c348 (.CLK(clknet_leaf_12_clk),
    .D(net13),
    .SCD(net850),
    .SCE(net157),
    .SET_B(clknet_1_0__leaf_net815),
    .Q(net284));
 sky130_fd_sc_hd__dfbbp_1 c349 (.CLK(clknet_leaf_12_clk),
    .D(net246),
    .RESET_B(clknet_1_0__leaf_net843),
    .SET_B(net157),
    .Q(net819),
    .Q_N(net285));
 sky130_fd_sc_hd__and3b_2 c350 (.A_N(clknet_1_1__leaf_net145),
    .B(net280),
    .C(net282),
    .X(net286));
 sky130_fd_sc_hd__or4bb_1 c351 (.A(net159),
    .B(net14),
    .C_N(net284),
    .D_N(net282),
    .X(net287));
 sky130_fd_sc_hd__or4bb_4 c352 (.A(net283),
    .B(net284),
    .C_N(net280),
    .D_N(net119),
    .X(net288));
 sky130_fd_sc_hd__or4bb_4 c353 (.A(clknet_1_0__leaf_net155),
    .B(net288),
    .C_N(net159),
    .D_N(net651),
    .X(net289));
 sky130_fd_sc_hd__mux4_2 c354 (.A0(net152),
    .A1(net288),
    .A2(clknet_1_1__leaf_net286),
    .A3(net40),
    .S0(net909),
    .S1(clknet_1_1__leaf_net289),
    .X(net290));
 sky130_fd_sc_hd__sdfxbp_1 c355 (.CLK(clknet_leaf_18_clk),
    .D(clknet_1_1__leaf_net228),
    .SCD(net290),
    .SCE(clknet_1_1__leaf_net145),
    .Q(net813),
    .Q_N(net291));
 sky130_fd_sc_hd__mux4_4 c356 (.A0(net284),
    .A1(net778),
    .A2(net281),
    .A3(net813),
    .S0(clknet_1_1__leaf_net269),
    .S1(clknet_1_1__leaf_net145),
    .X(net292));
 sky130_fd_sc_hd__mux4_2 c372 (.A0(net58),
    .A1(net284),
    .A2(clknet_1_1__leaf_net815),
    .A3(clknet_1_1__leaf_net843),
    .S0(net904),
    .S1(net847),
    .X(net835));
 sky130_fd_sc_hd__mux4_4 c373 (.A0(net747),
    .A1(net282),
    .A2(net176),
    .A3(clknet_1_0__leaf_net835),
    .S0(net824),
    .S1(net652),
    .X(net293));
 sky130_fd_sc_hd__mux4_2 c374 (.A0(net278),
    .A1(net8),
    .A2(net810),
    .A3(clknet_1_0__leaf_net812),
    .S0(net849),
    .S1(net653),
    .X(net294));
 sky130_fd_sc_hd__mux4_2 c375 (.A0(net782),
    .A1(clknet_1_1__leaf_net815),
    .A2(net282),
    .A3(clknet_1_0__leaf_net835),
    .S0(net651),
    .S1(net838),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net182),
    .A1(net830),
    .A2(net58),
    .A3(clknet_1_0__leaf_net835),
    .S0(net637),
    .S1(net836),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net287),
    .A1(net176),
    .A2(net182),
    .A3(clknet_1_0__leaf_net835),
    .S0(net891),
    .S1(net836),
    .X(net297));
 sky130_fd_sc_hd__nand2b_2 c378 (.A_N(net192),
    .B(net738),
    .Y(net298));
 sky130_fd_sc_hd__nand2b_1 c379 (.A_N(net189),
    .B(net200),
    .Y(net299));
 sky130_fd_sc_hd__dfrtn_1 c380 (.CLK_N(clknet_leaf_4_clk),
    .D(net793),
    .RESET_B(net299),
    .Q(net300));
 sky130_fd_sc_hd__dfrtp_4 c381 (.CLK(clknet_leaf_4_clk),
    .D(net299),
    .RESET_B(net187),
    .Q(net301));
 sky130_fd_sc_hd__and2_1 c382 (.A(net187),
    .B(net184),
    .X(net302));
 sky130_fd_sc_hd__nand2b_4 c383 (.A_N(net195),
    .B(net907),
    .Y(net303));
 sky130_fd_sc_hd__or3b_4 c384 (.A(net302),
    .B(net301),
    .C_N(net298),
    .X(net304));
 sky130_fd_sc_hd__and2b_2 c385 (.A_N(net185),
    .B(net890),
    .X(net305));
 sky130_fd_sc_hd__nand3b_1 c386 (.A_N(net304),
    .B(net298),
    .C(net305),
    .Y(net306));
 sky130_fd_sc_hd__nor2_1 c387 (.A(net184),
    .B(net305),
    .Y(net307));
 sky130_fd_sc_hd__or2b_2 c388 (.A(net305),
    .B_N(net306),
    .X(net308));
 sky130_fd_sc_hd__nand2b_1 c389 (.A_N(net306),
    .B(net889),
    .Y(net309));
 sky130_fd_sc_hd__nor3_2 c390 (.A(net194),
    .B(net877),
    .C(net303),
    .Y(net310));
 sky130_fd_sc_hd__or3_1 c391 (.A(net300),
    .B(net305),
    .C(net827),
    .X(net311));
 sky130_fd_sc_hd__a2111oi_1 c392 (.A1(net311),
    .A2(net883),
    .B1(net305),
    .C1(net304),
    .D1(net877),
    .Y(net312));
 sky130_fd_sc_hd__nor3b_1 c393 (.A(net869),
    .B(net889),
    .C_N(net305),
    .Y(net313));
 sky130_fd_sc_hd__sdfbbp_1 c394 (.CLK(clknet_leaf_4_clk),
    .D(net299),
    .RESET_B(net300),
    .SCD(net867),
    .SCE(net889),
    .SET_B(net308),
    .Q(net315),
    .Q_N(net314));
 sky130_fd_sc_hd__or3_4 c395 (.A(net200),
    .B(net307),
    .C(net867),
    .X(net316));
 sky130_fd_sc_hd__sdfstp_1 c396 (.CLK(clknet_leaf_4_clk),
    .D(net316),
    .SCD(net867),
    .SCE(net310),
    .SET_B(net918),
    .Q(net317));
 sky130_fd_sc_hd__sedfxbp_1 c397 (.CLK(clknet_leaf_4_clk),
    .D(net307),
    .DE(net317),
    .SCD(net298),
    .SCE(net316),
    .Q(net319),
    .Q_N(net318));
 sky130_fd_sc_hd__nand2b_2 c398 (.A_N(net313),
    .B(net201),
    .Y(net320));
 sky130_fd_sc_hd__or2b_1 c399 (.A(net756),
    .B_N(net68),
    .X(net321));
 sky130_fd_sc_hd__or4bb_1 c400 (.A(net759),
    .B(net212),
    .C_N(net202),
    .D_N(net221),
    .X(net322));
 sky130_fd_sc_hd__and2b_1 c401 (.A_N(net68),
    .B(net302),
    .X(net323));
 sky130_fd_sc_hd__and2_2 c402 (.A(net311),
    .B(net640),
    .X(net324));
 sky130_fd_sc_hd__or4bb_1 c403 (.A(net213),
    .B(net762),
    .C_N(net209),
    .D_N(net640),
    .X(net325));
 sky130_fd_sc_hd__and3b_4 c404 (.A_N(net322),
    .B(net307),
    .C(net883),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c405 (.A0(net748),
    .A1(net877),
    .A2(net325),
    .A3(net888),
    .S0(net324),
    .S1(net861),
    .X(net327));
 sky130_fd_sc_hd__nand3_1 c406 (.A(net323),
    .B(net220),
    .C(net861),
    .Y(net328));
 sky130_fd_sc_hd__a2111oi_1 c407 (.A1(net86),
    .A2(net213),
    .B1(net322),
    .C1(net861),
    .D1(net809),
    .Y(net329));
 sky130_fd_sc_hd__mux4_1 c408 (.A0(net328),
    .A1(net68),
    .A2(net221),
    .A3(net862),
    .S0(net756),
    .S1(net752),
    .X(net330));
 sky130_fd_sc_hd__a2111oi_1 c409 (.A1(net306),
    .A2(net327),
    .B1(net324),
    .C1(net861),
    .D1(net896),
    .Y(net331));
 sky130_fd_sc_hd__sdfxbp_1 c410 (.CLK(clknet_leaf_4_clk),
    .D(net330),
    .SCD(net861),
    .SCE(net311),
    .Q(net333),
    .Q_N(net332));
 sky130_fd_sc_hd__sedfxbp_1 c411 (.CLK(clknet_leaf_4_clk),
    .D(net948),
    .DE(net308),
    .SCD(net955),
    .SCE(net861),
    .Q(net335),
    .Q_N(net334));
 sky130_fd_sc_hd__or4bb_1 c412 (.A(net325),
    .B(net220),
    .C_N(net335),
    .D_N(net862),
    .X(net336));
 sky130_fd_sc_hd__sdfxtp_1 c413 (.CLK(clknet_leaf_3_clk),
    .D(net854),
    .SCD(net330),
    .SCE(net861),
    .Q(net337));
 sky130_fd_sc_hd__mux4_2 c414 (.A0(net335),
    .A1(net298),
    .A2(net221),
    .A3(net882),
    .S0(net862),
    .S1(net332),
    .X(net338));
 sky130_fd_sc_hd__a2111o_4 c415 (.A1(net956),
    .A2(net333),
    .B1(net322),
    .C1(net334),
    .D1(net861),
    .X(net339));
 sky130_fd_sc_hd__sdfxtp_1 c416 (.CLK(clknet_leaf_3_clk),
    .D(net330),
    .SCD(net927),
    .SCE(net861),
    .Q(net340));
 sky130_fd_sc_hd__sdfxtp_1 c417 (.CLK(clknet_leaf_3_clk),
    .D(net202),
    .SCD(net339),
    .SCE(net862),
    .Q(net341));
 sky130_fd_sc_hd__sedfxtp_4 c418 (.CLK(clknet_leaf_0_clk),
    .D(net213),
    .DE(net339),
    .SCD(net325),
    .SCE(net862),
    .Q(net342));
 sky130_fd_sc_hd__or3_4 c419 (.A(net338),
    .B(net342),
    .C(net861),
    .X(net343));
 sky130_fd_sc_hd__nand3_1 c420 (.A(net765),
    .B(net338),
    .C(net759),
    .Y(net344));
 sky130_fd_sc_hd__sedfxtp_1 c421 (.CLK(clknet_leaf_3_clk),
    .D(net866),
    .DE(net198),
    .SCD(net339),
    .SCE(net188),
    .Q(net345));
 sky130_fd_sc_hd__and3_2 c422 (.A(net321),
    .B(clknet_1_0__leaf_net236),
    .C(net646),
    .X(net817));
 sky130_fd_sc_hd__sedfxtp_1 c423 (.CLK(clknet_leaf_8_clk),
    .D(net941),
    .DE(net121),
    .SCD(net191),
    .SCE(net212),
    .Q(net346));
 sky130_fd_sc_hd__or4bb_1 c424 (.A(net336),
    .B(net206),
    .C_N(net739),
    .D_N(net782),
    .X(net347));
 sky130_fd_sc_hd__o2111ai_1 c425 (.A1(net341),
    .A2(net765),
    .B1(net782),
    .C1(net234),
    .D1(net862),
    .Y(net348));
 sky130_fd_sc_hd__or3b_1 c426 (.A(net327),
    .B(net321),
    .C_N(net782),
    .X(net349));
 sky130_fd_sc_hd__or3b_1 c427 (.A(net919),
    .B(net336),
    .C_N(net863),
    .X(net350));
 sky130_fd_sc_hd__mux4_2 c428 (.A0(net98),
    .A1(net227),
    .A2(net321),
    .A3(net866),
    .S0(net220),
    .S1(net303),
    .X(net351));
 sky130_fd_sc_hd__sdfbbn_1 c429 (.CLK_N(clknet_leaf_9_clk),
    .D(net349),
    .RESET_B(net212),
    .SCD(clknet_1_0__leaf_net240),
    .SCE(net790),
    .SET_B(net892),
    .Q(net353),
    .Q_N(net352));
 sky130_fd_sc_hd__dfbbn_1 c430 (.CLK_N(clknet_leaf_3_clk),
    .D(net350),
    .RESET_B(net128),
    .SET_B(net323),
    .Q(net355),
    .Q_N(net354));
 sky130_fd_sc_hd__sdfrbp_1 c431 (.CLK(clknet_leaf_3_clk),
    .D(net348),
    .RESET_B(net198),
    .SCD(net350),
    .SCE(net352),
    .Q(net357),
    .Q_N(net356));
 sky130_fd_sc_hd__sdfbbn_1 c432 (.CLK_N(clknet_leaf_9_clk),
    .D(net937),
    .RESET_B(net234),
    .SCD(net356),
    .SCE(clknet_1_1__leaf_net238),
    .SET_B(net939),
    .Q(net359),
    .Q_N(net358));
 sky130_fd_sc_hd__sdfbbp_1 c433 (.CLK(clknet_leaf_3_clk),
    .D(net929),
    .RESET_B(net756),
    .SCD(net347),
    .SCE(net354),
    .SET_B(net350),
    .Q(net361),
    .Q_N(net360));
 sky130_fd_sc_hd__or4bb_1 c434 (.A(net337),
    .B(net355),
    .C_N(net360),
    .D_N(net866),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net298),
    .A1(net357),
    .A2(net353),
    .A3(net765),
    .S0(net119),
    .S1(net878),
    .X(net837));
 sky130_fd_sc_hd__sdfrbp_2 c436 (.CLK(clknet_leaf_2_clk),
    .D(net344),
    .RESET_B(net917),
    .SCD(net355),
    .SCE(net872),
    .Q(net364),
    .Q_N(net363));
 sky130_fd_sc_hd__a2111o_4 c437 (.A1(net355),
    .A2(net364),
    .B1(net352),
    .C1(net872),
    .D1(net883),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net364),
    .A1(net346),
    .A2(net356),
    .A3(net354),
    .S0(net365),
    .S1(net872),
    .X(net366));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net227),
    .A1(net873),
    .A2(net366),
    .A3(net317),
    .S0(net356),
    .S1(net354),
    .X(net367));
 sky130_fd_sc_hd__mux4_2 c440 (.A0(net347),
    .A1(net366),
    .A2(net357),
    .A3(net351),
    .S0(net310),
    .S1(net363),
    .X(net368));
 sky130_fd_sc_hd__and2_1 c441 (.A(net353),
    .B(net905),
    .X(net369));
 sky130_fd_sc_hd__or2b_2 c442 (.A(net359),
    .B_N(net746),
    .X(net370));
 sky130_fd_sc_hd__nand3_2 c443 (.A(clknet_1_0__leaf_net255),
    .B(net863),
    .C(net873),
    .Y(net371));
 sky130_fd_sc_hd__sdfbbn_1 c444 (.CLK_N(clknet_leaf_9_clk),
    .D(net361),
    .RESET_B(net364),
    .SCD(net256),
    .SCE(net358),
    .SET_B(net339),
    .Q(net372));
 sky130_fd_sc_hd__or2b_2 c445 (.A(net372),
    .B_N(net886),
    .X(net373));
 sky130_fd_sc_hd__nand3b_4 c446 (.A_N(net369),
    .B(net868),
    .C(net873),
    .Y(net823));
 sky130_fd_sc_hd__nand3_1 c447 (.A(net373),
    .B(net205),
    .C(net886),
    .Y(net374));
 sky130_fd_sc_hd__o2111ai_4 c448 (.A1(net373),
    .A2(net364),
    .B1(net886),
    .C1(net247),
    .D1(net873),
    .Y(net375));
 sky130_fd_sc_hd__and3b_1 c449 (.A_N(net371),
    .B(net964),
    .C(net375),
    .X(net376));
 sky130_fd_sc_hd__nand2b_1 c450 (.A_N(net375),
    .B(net363),
    .Y(net377));
 sky130_fd_sc_hd__or4bb_1 c451 (.A(net302),
    .B(clknet_1_0__leaf_net255),
    .C_N(net373),
    .D_N(net886),
    .X(net378));
 sky130_fd_sc_hd__nand3_4 c452 (.A(net248),
    .B(net886),
    .C(clknet_1_0__leaf_net378),
    .Y(net379));
 sky130_fd_sc_hd__mux4_2 c453 (.A0(clknet_1_0__leaf_net378),
    .A1(net784),
    .A2(net373),
    .A3(net375),
    .S0(net905),
    .S1(net873),
    .X(net380));
 sky130_fd_sc_hd__or3_1 c454 (.A(net377),
    .B(net18),
    .C(clknet_1_0__leaf_net378),
    .X(net381));
 sky130_fd_sc_hd__mux4_4 c455 (.A0(net376),
    .A1(clknet_1_0__leaf_net261),
    .A2(net18),
    .A3(net375),
    .S0(clknet_1_1__leaf_net378),
    .S1(net892),
    .X(net382));
 sky130_fd_sc_hd__mux4_2 c456 (.A0(net374),
    .A1(clknet_1_0__leaf_net378),
    .A2(net363),
    .A3(clknet_1_1__leaf_net379),
    .S0(clknet_1_0__leaf_net381),
    .S1(net892),
    .X(net383));
 sky130_fd_sc_hd__sdfbbn_2 c457 (.CLK_N(clknet_leaf_19_clk),
    .D(clknet_1_0__leaf_net261),
    .RESET_B(clknet_1_1__leaf_net378),
    .SCD(net905),
    .SCE(net377),
    .SET_B(net656),
    .Q(net385),
    .Q_N(net384));
 sky130_fd_sc_hd__mux4_2 c458 (.A0(clknet_1_1__leaf_net381),
    .A1(net375),
    .A2(clknet_1_0__leaf_net269),
    .A3(net18),
    .S0(net886),
    .S1(net646),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net898),
    .A1(clknet_1_1__leaf_net378),
    .A2(net384),
    .A3(net343),
    .S0(net375),
    .S1(net656),
    .X(net387));
 sky130_fd_sc_hd__o2111ai_1 c460 (.A1(net353),
    .A2(net367),
    .B1(net873),
    .C1(net654),
    .D1(net655),
    .Y(net388));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net388),
    .A1(net339),
    .A2(clknet_1_1__leaf_net378),
    .A3(clknet_1_1__leaf_net238),
    .S0(net384),
    .S1(net655),
    .X(net389));
 sky130_fd_sc_hd__nor3b_2 c462 (.A(net362),
    .B(clknet_1_0__leaf_net818),
    .C_N(net832),
    .Y(net801));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(clknet_1_0__leaf_net269),
    .A1(net163),
    .A2(net127),
    .A3(clknet_1_0__leaf_net823),
    .S0(net733),
    .S1(clknet_1_0__leaf_net815),
    .X(net390));
 sky130_fd_sc_hd__mux4_2 c464 (.A0(net36),
    .A1(clknet_1_0__leaf_net818),
    .A2(net886),
    .A3(clknet_1_0__leaf_net815),
    .S0(clknet_1_1__leaf_net379),
    .S1(net660),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net279),
    .A1(clknet_1_1__leaf_net238),
    .A2(clknet_1_0__leaf_net801),
    .A3(clknet_1_1__leaf_net289),
    .S0(net903),
    .S1(net657),
    .X(net392));
 sky130_fd_sc_hd__sdfbbp_1 c466 (.CLK(clknet_leaf_19_clk),
    .D(net942),
    .RESET_B(clknet_1_0__leaf_net801),
    .SCD(net931),
    .SCE(net661),
    .SET_B(net663),
    .Q(net393));
 sky130_fd_sc_hd__and3b_1 c467 (.A_N(net206),
    .B(clknet_1_0__leaf_net829),
    .C(net964),
    .X(net394));
 sky130_fd_sc_hd__and3b_2 c468 (.A_N(net271),
    .B(net882),
    .C(net663),
    .X(net395));
 sky130_fd_sc_hd__nand3b_1 c469 (.A_N(net270),
    .B(net662),
    .C(net663),
    .Y(net396));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net367),
    .A1(clknet_1_0__leaf_net829),
    .A2(net864),
    .A3(net291),
    .S0(net395),
    .S1(net832),
    .X(net852));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net396),
    .A1(net274),
    .A2(net304),
    .A3(net395),
    .S0(net370),
    .S1(net270),
    .X(net397));
 sky130_fd_sc_hd__and3_1 c472 (.A(net395),
    .B(net304),
    .C(net658),
    .X(net833));
 sky130_fd_sc_hd__and3_4 c473 (.A(net274),
    .B(net291),
    .C(net658),
    .X(net398));
 sky130_fd_sc_hd__and3b_2 c474 (.A_N(net317),
    .B(net36),
    .C(net868),
    .X(net807));
 sky130_fd_sc_hd__and3b_1 c475 (.A_N(net36),
    .B(net303),
    .C(net395),
    .X(net399));
 sky130_fd_sc_hd__mux4_4 c476 (.A0(net303),
    .A1(net395),
    .A2(net863),
    .A3(net398),
    .S0(clknet_1_0__leaf_net801),
    .S1(net832),
    .X(net400));
 sky130_fd_sc_hd__nor3b_1 c477 (.A(net393),
    .B(net807),
    .C_N(net813),
    .Y(net401));
 sky130_fd_sc_hd__mux4_2 c478 (.A0(net399),
    .A1(net965),
    .A2(net881),
    .A3(clknet_1_0__leaf_net852),
    .S0(net882),
    .S1(net661),
    .X(net402));
 sky130_fd_sc_hd__mux4_2 c479 (.A0(net401),
    .A1(clknet_1_0__leaf_net286),
    .A2(net395),
    .A3(net279),
    .S0(net398),
    .S1(net663),
    .X(net403));
 sky130_fd_sc_hd__mux4_4 c480 (.A0(net397),
    .A1(net873),
    .A2(net395),
    .A3(clknet_1_0__leaf_net852),
    .S0(clknet_1_1__leaf_net801),
    .S1(net665),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net778),
    .A1(clknet_1_0__leaf_net823),
    .A2(net395),
    .A3(clknet_1_1__leaf_net801),
    .S0(net667),
    .S1(net828),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net395),
    .A1(clknet_1_1__leaf_net815),
    .A2(net36),
    .A3(net881),
    .S0(net828),
    .S1(net668),
    .X(net406));
 sky130_fd_sc_hd__and2b_1 c504 (.A_N(net300),
    .B(net953),
    .X(net407));
 sky130_fd_sc_hd__inv_1 c505 (.A(net922),
    .Y(net408));
 sky130_fd_sc_hd__nand2b_2 c506 (.A_N(net732),
    .B(net408),
    .Y(net409));
 sky130_fd_sc_hd__nand2b_2 c507 (.A_N(net312),
    .B(net907),
    .Y(net410));
 sky130_fd_sc_hd__dfbbn_2 c508 (.CLK_N(clknet_leaf_32_clk),
    .D(net316),
    .RESET_B(net410),
    .SET_B(net408),
    .Q(net412),
    .Q_N(net411));
 sky130_fd_sc_hd__nor2b_2 c509 (.A(net309),
    .B_N(net412),
    .Y(net413));
 sky130_fd_sc_hd__clkbuf_2 c510 (.A(net922),
    .X(net414));
 sky130_fd_sc_hd__a2111o_1 c511 (.A1(net407),
    .A2(net408),
    .B1(net413),
    .C1(net414),
    .D1(net410),
    .X(net415));
 sky130_fd_sc_hd__or2b_1 c512 (.A(net412),
    .B_N(net408),
    .X(net416));
 sky130_fd_sc_hd__nand3b_4 c513 (.A_N(net201),
    .B(net414),
    .C(net883),
    .Y(net417));
 sky130_fd_sc_hd__and2b_1 c514 (.A_N(net410),
    .B(net315),
    .X(net418));
 sky130_fd_sc_hd__nor3_1 c515 (.A(net416),
    .B(net308),
    .C(net415),
    .Y(net419));
 sky130_fd_sc_hd__dfrtp_4 c516 (.CLK(clknet_leaf_30_clk),
    .D(net419),
    .RESET_B(net415),
    .Q(net420));
 sky130_fd_sc_hd__nor3_1 c517 (.A(net409),
    .B(net418),
    .C(net414),
    .Y(net421));
 sky130_fd_sc_hd__nor2b_1 c518 (.A(net421),
    .B_N(net414),
    .Y(net422));
 sky130_fd_sc_hd__dfbbp_1 c519 (.CLK(clknet_leaf_32_clk),
    .D(net407),
    .RESET_B(net421),
    .SET_B(net316),
    .Q(net424),
    .Q_N(net423));
 sky130_fd_sc_hd__sdfxbp_1 c520 (.CLK(clknet_leaf_30_clk),
    .D(net419),
    .SCD(net422),
    .SCE(net423),
    .Q(net426),
    .Q_N(net425));
 sky130_fd_sc_hd__mux4_1 c521 (.A0(net426),
    .A1(net859),
    .A2(net309),
    .A3(net411),
    .S0(net308),
    .S1(net316),
    .X(net427));
 sky130_fd_sc_hd__sdfxbp_1 c522 (.CLK(clknet_leaf_31_clk),
    .D(net422),
    .SCD(net424),
    .SCE(net415),
    .Q(net429),
    .Q_N(net428));
 sky130_fd_sc_hd__mux4_2 c523 (.A0(net914),
    .A1(net413),
    .A2(net859),
    .A3(net414),
    .S0(net893),
    .S1(net952),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(net421),
    .A1(net428),
    .A2(net417),
    .A3(net316),
    .S0(net409),
    .S1(net669),
    .X(net431));
 sky130_fd_sc_hd__nand3b_1 c525 (.A_N(net408),
    .B(net883),
    .C(net413),
    .Y(net432));
 sky130_fd_sc_hd__and3_1 c526 (.A(net738),
    .B(net220),
    .C(net432),
    .X(net433));
 sky130_fd_sc_hd__sdfxtp_1 c527 (.CLK(clknet_leaf_32_clk),
    .D(net414),
    .SCD(net308),
    .SCE(net430),
    .Q(net434));
 sky130_fd_sc_hd__and3_1 c528 (.A(net429),
    .B(net325),
    .C(net434),
    .X(net435));
 sky130_fd_sc_hd__dfrtp_4 c529 (.CLK(clknet_leaf_32_clk),
    .D(net768),
    .RESET_B(net430),
    .Q(net436));
 sky130_fd_sc_hd__dfsbp_1 c530 (.CLK(clknet_leaf_0_clk),
    .D(net308),
    .SET_B(net320),
    .Q(net438),
    .Q_N(net437));
 sky130_fd_sc_hd__and3b_1 c531 (.A_N(net432),
    .B(net436),
    .C(clknet_1_1__leaf_net670),
    .X(net439));
 sky130_fd_sc_hd__sdfxtp_1 c532 (.CLK(clknet_leaf_0_clk),
    .D(net888),
    .SCD(net936),
    .SCE(net343),
    .Q(net440));
 sky130_fd_sc_hd__nor3b_1 c533 (.A(net896),
    .B(net436),
    .C_N(net888),
    .Y(net441));
 sky130_fd_sc_hd__sdfxtp_1 c534 (.CLK(clknet_leaf_31_clk),
    .D(net441),
    .SCD(clknet_1_0__leaf_net439),
    .SCE(net949),
    .Q(net442));
 sky130_fd_sc_hd__dfbbn_1 c535 (.CLK_N(clknet_leaf_31_clk),
    .D(net436),
    .RESET_B(net442),
    .SET_B(clknet_1_0__leaf_net439),
    .Q(net444),
    .Q_N(net443));
 sky130_fd_sc_hd__dfbbn_1 c536 (.CLK_N(clknet_leaf_32_clk),
    .D(net430),
    .RESET_B(net441),
    .SET_B(net436),
    .Q(net445));
 sky130_fd_sc_hd__or3b_2 c537 (.A(net435),
    .B(net436),
    .C_N(net870),
    .X(net446));
 sky130_fd_sc_hd__o2111a_1 c538 (.A1(net445),
    .A2(net442),
    .B1(net443),
    .C1(net436),
    .D1(net446),
    .X(net447));
 sky130_fd_sc_hd__o2111a_4 c539 (.A1(net324),
    .A2(net870),
    .B1(net440),
    .C1(net446),
    .D1(net188),
    .X(net448));
 sky130_fd_sc_hd__dfbbp_1 c540 (.CLK(clknet_leaf_0_clk),
    .D(net433),
    .RESET_B(net446),
    .SET_B(net444),
    .Q(net450),
    .Q_N(net449));
 sky130_fd_sc_hd__sdfbbn_2 c541 (.CLK_N(clknet_leaf_0_clk),
    .D(net305),
    .RESET_B(net436),
    .SCD(net448),
    .SCE(clknet_1_1__leaf_net439),
    .SET_B(net434),
    .Q(net452),
    .Q_N(net451));
 sky130_fd_sc_hd__a2111oi_4 c542 (.A1(net447),
    .A2(net324),
    .B1(net450),
    .C1(net888),
    .D1(net451),
    .Y(net799));
 sky130_fd_sc_hd__a2111o_1 c543 (.A1(net198),
    .A2(net452),
    .B1(net324),
    .C1(net858),
    .D1(net446),
    .X(net453));
 sky130_fd_sc_hd__sdfbbn_1 c544 (.CLK_N(clknet_leaf_31_clk),
    .D(net442),
    .RESET_B(net799),
    .SCD(net452),
    .SCE(net450),
    .SET_B(net453),
    .Q(net454));
 sky130_fd_sc_hd__sdfbbp_1 c545 (.CLK(clknet_leaf_0_clk),
    .D(net454),
    .RESET_B(net453),
    .SCD(net339),
    .SCE(net438),
    .SET_B(net451),
    .Q(net456),
    .Q_N(net455));
 sky130_fd_sc_hd__sdfxbp_1 c546 (.CLK(clknet_leaf_0_clk),
    .D(net947),
    .SCD(net343),
    .SCE(net878),
    .Q(net458),
    .Q_N(net457));
 sky130_fd_sc_hd__and3b_2 c547 (.A_N(net778),
    .B(net365),
    .C(net752),
    .X(net459));
 sky130_fd_sc_hd__sdfbbn_1 c548 (.CLK_N(clknet_leaf_1_clk),
    .D(net458),
    .RESET_B(net870),
    .SCD(net417),
    .SCE(net459),
    .SET_B(net440),
    .Q(net461),
    .Q_N(net460));
 sky130_fd_sc_hd__or3_1 c549 (.A(net461),
    .B(net452),
    .C(net434),
    .X(net462));
 sky130_fd_sc_hd__mux4_2 c550 (.A0(clknet_1_0__leaf_net240),
    .A1(net462),
    .A2(net434),
    .A3(net451),
    .S0(net857),
    .S1(net878),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(net440),
    .A1(net351),
    .A2(net338),
    .A3(net449),
    .S0(net459),
    .S1(net339),
    .X(net464));
 sky130_fd_sc_hd__a2111oi_1 c552 (.A1(net234),
    .A2(net858),
    .B1(net459),
    .C1(net437),
    .D1(net460),
    .Y(net465));
 sky130_fd_sc_hd__sdfbbn_1 c553 (.CLK_N(clknet_leaf_1_clk),
    .D(net954),
    .RESET_B(net412),
    .SCD(net933),
    .SCE(net314),
    .SET_B(clknet_1_0__leaf_net671),
    .Q(net467),
    .Q_N(net466));
 sky130_fd_sc_hd__sdfbbp_1 c554 (.CLK(clknet_leaf_1_clk),
    .D(net221),
    .RESET_B(net878),
    .SCD(net351),
    .SCE(net853),
    .SET_B(clknet_1_0__leaf_net671),
    .Q(net468));
 sky130_fd_sc_hd__sdfbbn_1 c555 (.CLK_N(clknet_leaf_1_clk),
    .D(net752),
    .RESET_B(net878),
    .SCD(net944),
    .SCE(net954),
    .SET_B(clknet_1_0__leaf_net671),
    .Q(net470),
    .Q_N(net469));
 sky130_fd_sc_hd__sdfxbp_2 c556 (.CLK(clknet_leaf_2_clk),
    .D(net467),
    .SCD(net417),
    .SCE(net342),
    .Q(net804),
    .Q_N(net471));
 sky130_fd_sc_hd__o2111a_1 c557 (.A1(net459),
    .A2(net434),
    .B1(net804),
    .C1(net469),
    .D1(net873),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net470),
    .A1(net365),
    .A2(net954),
    .A3(net412),
    .S0(clknet_1_1__leaf_net463),
    .S1(net471),
    .X(net473));
 sky130_fd_sc_hd__mux4_4 c559 (.A0(net472),
    .A1(net870),
    .A2(net732),
    .A3(net669),
    .S0(clknet_1_0__leaf_net671),
    .S1(clknet_1_1__leaf_net672),
    .X(net474));
 sky130_fd_sc_hd__mux4_2 c560 (.A0(net883),
    .A1(clknet_1_0__leaf_net474),
    .A2(net853),
    .A3(net457),
    .S0(net669),
    .S1(clknet_1_1__leaf_net672),
    .X(net475));
 sky130_fd_sc_hd__a2111oi_4 c561 (.A1(net468),
    .A2(net804),
    .B1(net450),
    .C1(clknet_1_1__leaf_net672),
    .D1(clknet_1_0__leaf_net474),
    .Y(net476));
 sky130_fd_sc_hd__mux4_4 c562 (.A0(clknet_1_1__leaf_net474),
    .A1(net338),
    .A2(net459),
    .A3(net471),
    .S0(clknet_1_0__leaf_net476),
    .S1(clknet_1_1__leaf_net672),
    .X(net477));
 sky130_fd_sc_hd__mux4_4 c563 (.A0(clknet_1_0__leaf_net476),
    .A1(net459),
    .A2(clknet_1_1__leaf_net474),
    .A3(net351),
    .S0(net471),
    .S1(net675),
    .X(net478));
 sky130_fd_sc_hd__mux4_4 c564 (.A0(net315),
    .A1(net338),
    .A2(net411),
    .A3(clknet_1_0__leaf_net474),
    .S0(net673),
    .S1(net674),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(clknet_1_0__leaf_net479),
    .A1(net472),
    .A2(net804),
    .A3(clknet_1_1__leaf_net474),
    .S0(net853),
    .S1(net675),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net865),
    .A1(clknet_1_1__leaf_net479),
    .A2(net784),
    .A3(net674),
    .S0(net677),
    .S1(net678),
    .X(net481));
 sky130_fd_sc_hd__sdfbbn_2 c567 (.CLK_N(clknet_leaf_25_clk),
    .D(net351),
    .RESET_B(net926),
    .SCD(net265),
    .SCE(net893),
    .SET_B(net339),
    .Q(net483),
    .Q_N(net482));
 sky130_fd_sc_hd__or3b_1 c568 (.A(net18),
    .B(net804),
    .C_N(net892),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net484),
    .A1(net385),
    .A2(net795),
    .A3(net18),
    .S0(net443),
    .S1(net856),
    .X(net485));
 sky130_fd_sc_hd__sdfbbp_1 c570 (.CLK(clknet_leaf_25_clk),
    .D(net265),
    .RESET_B(net343),
    .SCD(clknet_1_0__leaf_net142),
    .SCE(net339),
    .SET_B(net872),
    .Q(net487),
    .Q_N(net486));
 sky130_fd_sc_hd__mux4_4 c571 (.A0(net339),
    .A1(net448),
    .A2(net119),
    .A3(clknet_1_0__leaf_net142),
    .S0(clknet_1_1__leaf_net379),
    .S1(net482),
    .X(net488));
 sky130_fd_sc_hd__mux4_2 c572 (.A0(net484),
    .A1(clknet_1_0__leaf_net142),
    .A2(net370),
    .A3(net448),
    .S0(net676),
    .S1(net680),
    .X(net489));
 sky130_fd_sc_hd__nor3b_2 c573 (.A(net265),
    .B(net677),
    .C_N(net680),
    .Y(net490));
 sky130_fd_sc_hd__mux4_4 c574 (.A0(net487),
    .A1(net256),
    .A2(net455),
    .A3(clknet_1_0__leaf_net489),
    .S0(net870),
    .S1(net872),
    .X(net491));
 sky130_fd_sc_hd__a2111o_1 c575 (.A1(net342),
    .A2(net486),
    .B1(net490),
    .C1(net872),
    .D1(net448),
    .X(net492));
 sky130_fd_sc_hd__or4bb_1 c576 (.A(net490),
    .B(net342),
    .C_N(net492),
    .D_N(net873),
    .X(net493));
 sky130_fd_sc_hd__sdfxtp_1 c577 (.CLK(clknet_leaf_25_clk),
    .D(net485),
    .SCD(net351),
    .SCE(net448),
    .Q(net494));
 sky130_fd_sc_hd__mux4_4 c578 (.A0(net212),
    .A1(net343),
    .A2(net494),
    .A3(net482),
    .S0(net455),
    .S1(clknet_1_1__leaf_net476),
    .X(net495));
 sky130_fd_sc_hd__or4bb_2 c579 (.A(net494),
    .B(net448),
    .C_N(net897),
    .D_N(net326),
    .X(net496));
 sky130_fd_sc_hd__mux4_4 c580 (.A0(net493),
    .A1(net492),
    .A2(net264),
    .A3(net384),
    .S0(clknet_1_0__leaf_net142),
    .S1(net679),
    .X(net497));
 sky130_fd_sc_hd__or3_1 c581 (.A(net492),
    .B(net868),
    .C(net342),
    .X(net498));
 sky130_fd_sc_hd__mux4_4 c582 (.A0(clknet_1_0__leaf_net491),
    .A1(net856),
    .A2(net492),
    .A3(net351),
    .S0(net483),
    .S1(net493),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net380),
    .A1(net739),
    .A2(clknet_1_1__leaf_net491),
    .A3(net496),
    .S0(net448),
    .S1(clknet_1_0__leaf_net142),
    .X(net500));
 sky130_fd_sc_hd__mux4_4 c584 (.A0(net448),
    .A1(clknet_1_0__leaf_net142),
    .A2(net471),
    .A3(net84),
    .S0(net683),
    .S1(net686),
    .X(net501));
 sky130_fd_sc_hd__mux4_2 c585 (.A0(net498),
    .A1(clknet_1_0__leaf_net501),
    .A2(net893),
    .A3(clknet_1_1__leaf_net379),
    .S0(net492),
    .S1(net683),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(clknet_1_1__leaf_net501),
    .A1(clknet_1_0__leaf_net142),
    .A2(net892),
    .A3(net891),
    .S0(net680),
    .S1(net685),
    .X(net503));
 sky130_fd_sc_hd__mux4_2 c587 (.A0(net264),
    .A1(net891),
    .A2(net679),
    .A3(net680),
    .S0(net681),
    .S1(net687),
    .X(net504));
 sky130_fd_sc_hd__mux4_4 c588 (.A0(net893),
    .A1(net385),
    .A2(net490),
    .A3(net288),
    .S0(net874),
    .S1(net684),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net505),
    .A1(net398),
    .A2(clknet_1_1__leaf_net289),
    .A3(net385),
    .S0(net881),
    .S1(clknet_1_0__leaf_net394),
    .X(net506));
 sky130_fd_sc_hd__mux4_2 c590 (.A0(clknet_1_1__leaf_net394),
    .A1(net881),
    .A2(net964),
    .A3(net504),
    .S0(clknet_1_0__leaf_net801),
    .S1(net482),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net448),
    .A1(net412),
    .A2(net163),
    .A3(net881),
    .S0(net504),
    .S1(net863),
    .X(net508));
 sky130_fd_sc_hd__mux4_2 c592 (.A0(net490),
    .A1(clknet_1_0__leaf_net379),
    .A2(net863),
    .A3(clknet_1_0__leaf_net801),
    .S0(net679),
    .S1(net688),
    .X(net509));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net462),
    .A1(net506),
    .A2(clknet_1_0__leaf_net394),
    .A3(net163),
    .S0(net288),
    .S1(clknet_1_1__leaf_net476),
    .X(net510));
 sky130_fd_sc_hd__mux4_2 c594 (.A0(net790),
    .A1(net868),
    .A2(net412),
    .A3(net881),
    .S0(net807),
    .S1(net681),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net882),
    .A1(net504),
    .A2(net897),
    .A3(net664),
    .S0(net687),
    .S1(net688),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net870),
    .A1(net865),
    .A2(clknet_1_0__leaf_net289),
    .A3(net304),
    .S0(net688),
    .S1(clknet_1_0__leaf_net689),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net406),
    .A1(net886),
    .A2(net398),
    .A3(net304),
    .S0(net664),
    .S1(net666),
    .X(net514));
 sky130_fd_sc_hd__mux4_4 c598 (.A0(net512),
    .A1(net882),
    .A2(clknet_1_1__leaf_net514),
    .A3(clknet_1_1__leaf_net289),
    .S0(net891),
    .S1(net684),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(clknet_1_0__leaf_net514),
    .A1(net398),
    .A2(net881),
    .A3(net163),
    .S0(net886),
    .S1(net411),
    .X(net516));
 sky130_fd_sc_hd__mux4_4 c600 (.A0(net964),
    .A1(net288),
    .A2(clknet_1_0__leaf_net289),
    .A3(net511),
    .S0(net482),
    .S1(clknet_1_0__leaf_net690),
    .X(net517));
 sky130_fd_sc_hd__mux4_2 c601 (.A0(net163),
    .A1(net288),
    .A2(net398),
    .A3(net856),
    .S0(net882),
    .S1(net688),
    .X(net811));
 sky130_fd_sc_hd__mux4_2 c602 (.A0(net868),
    .A1(net511),
    .A2(net163),
    .A3(clknet_1_0__leaf_net801),
    .S0(net966),
    .S1(net681),
    .X(net518));
 sky130_fd_sc_hd__mux4_2 c603 (.A0(clknet_1_1__leaf_net801),
    .A1(net411),
    .A2(net892),
    .A3(clknet_1_1__leaf_net690),
    .S0(clknet_1_1__leaf_net691),
    .S1(net693),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net220),
    .A1(net790),
    .A2(clknet_1_1__leaf_net513),
    .A3(net684),
    .S0(clknet_1_0__leaf_net689),
    .S1(net694),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net517),
    .A1(net504),
    .A2(clknet_1_0__leaf_net514),
    .A3(net865),
    .S0(net694),
    .S1(net695),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net452),
    .A1(net119),
    .A2(net891),
    .A3(net687),
    .S0(net688),
    .S1(net692),
    .X(net522));
 sky130_fd_sc_hd__mux4_2 c607 (.A0(net119),
    .A1(clknet_1_1__leaf_net852),
    .A2(clknet_1_1__leaf_net513),
    .A3(net511),
    .S0(net897),
    .S1(net696),
    .X(net523));
 sky130_fd_sc_hd__mux4_4 c608 (.A0(net522),
    .A1(net411),
    .A2(net688),
    .A3(clknet_1_1__leaf_net689),
    .S0(net797),
    .S1(net698),
    .X(net808));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net771),
    .A1(net781),
    .A2(net785),
    .A3(net788),
    .S0(net763),
    .S1(net782),
    .X(net0));
 sky130_fd_sc_hd__nor2b_1 c63 (.A(net775),
    .B_N(net3),
    .Y(net1));
 sky130_fd_sc_hd__or2_1 c630 (.A(net907),
    .B(net409),
    .X(net524));
 sky130_fd_sc_hd__and2_2 c631 (.A(net416),
    .B(net69),
    .X(net525));
 sky130_fd_sc_hd__and3b_2 c632 (.A_N(net186),
    .B(net409),
    .C(net524),
    .X(net526));
 sky130_fd_sc_hd__and2b_2 c633 (.A_N(net424),
    .B(net410),
    .X(net826));
 sky130_fd_sc_hd__nor3b_1 c634 (.A(net526),
    .B(net409),
    .C_N(net860),
    .Y(net527));
 sky130_fd_sc_hd__or4bb_2 c635 (.A(net410),
    .B(net525),
    .C_N(net186),
    .D_N(net860),
    .X(net528));
 sky130_fd_sc_hd__and3_1 c636 (.A(net525),
    .B(net425),
    .C(net860),
    .X(net529));
 sky130_fd_sc_hd__or4bb_1 c637 (.A(net529),
    .B(net528),
    .C_N(net413),
    .D_N(clknet_1_0__leaf_net670),
    .X(net530));
 sky130_fd_sc_hd__and3_1 c638 (.A(net524),
    .B(net186),
    .C(net525),
    .X(net531));
 sky130_fd_sc_hd__or4bb_1 c639 (.A(net531),
    .B(net525),
    .C_N(net527),
    .D_N(net409),
    .X(net532));
 sky130_fd_sc_hd__nand2_2 c64 (.A(net774),
    .B(net782),
    .Y(net2));
 sky130_fd_sc_hd__nor3_1 c640 (.A(net528),
    .B(net301),
    .C(net896),
    .Y(net533));
 sky130_fd_sc_hd__dfsbp_1 c641 (.CLK(clknet_leaf_29_clk),
    .D(net532),
    .SET_B(net528),
    .Q(net535),
    .Q_N(net534));
 sky130_fd_sc_hd__sdfxtp_1 c642 (.CLK(clknet_leaf_30_clk),
    .D(net415),
    .SCD(net531),
    .SCE(clknet_1_0__leaf_net530),
    .Q(net536));
 sky130_fd_sc_hd__nor2b_1 c643 (.A(net426),
    .B_N(net855),
    .Y(net537));
 sky130_fd_sc_hd__sdfrtn_1 c644 (.CLK_N(clknet_leaf_29_clk),
    .D(net533),
    .RESET_B(net535),
    .SCD(net855),
    .SCE(net906),
    .Q(net538));
 sky130_fd_sc_hd__sdfxtp_2 c645 (.CLK(clknet_leaf_30_clk),
    .D(net418),
    .SCD(clknet_1_0__leaf_net530),
    .SCE(net860),
    .Q(net539));
 sky130_fd_sc_hd__dfbbn_1 c646 (.CLK_N(clknet_leaf_29_clk),
    .D(net537),
    .RESET_B(net533),
    .SET_B(net526),
    .Q(net541),
    .Q_N(net540));
 sky130_fd_sc_hd__sdfrtp_1 c647 (.CLK(clknet_leaf_29_clk),
    .D(net532),
    .RESET_B(net538),
    .SCD(net536),
    .SCE(net524),
    .Q(net542));
 sky130_fd_sc_hd__mux4_2 c648 (.A0(net542),
    .A1(net527),
    .A2(net540),
    .A3(net410),
    .S0(net534),
    .S1(net524),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net541),
    .A1(net536),
    .A2(net537),
    .A3(net301),
    .S0(net543),
    .S1(net539),
    .X(net544));
 sky130_fd_sc_hd__or3_4 c65 (.A(net764),
    .B(net755),
    .C(net790),
    .X(net3));
 sky130_fd_sc_hd__mux4_1 c650 (.A0(net538),
    .A1(net524),
    .A2(net542),
    .A3(net543),
    .S0(net410),
    .S1(net531),
    .X(net545));
 sky130_fd_sc_hd__sdfrtp_1 c651 (.CLK(clknet_leaf_31_clk),
    .D(net209),
    .RESET_B(net528),
    .SCD(net417),
    .SCE(net893),
    .Q(net546));
 sky130_fd_sc_hd__or3b_2 c652 (.A(net340),
    .B(net449),
    .C_N(clknet_1_0__leaf_net670),
    .X(net547));
 sky130_fd_sc_hd__nand2b_1 c653 (.A_N(net340),
    .B(net536),
    .Y(net548));
 sky130_fd_sc_hd__dfbbn_1 c654 (.CLK_N(clknet_leaf_30_clk),
    .D(net320),
    .RESET_B(net221),
    .SET_B(net699),
    .Q(net550),
    .Q_N(net549));
 sky130_fd_sc_hd__dfbbp_1 c655 (.CLK(clknet_leaf_29_clk),
    .D(net413),
    .RESET_B(net526),
    .SET_B(net543),
    .Q(net551));
 sky130_fd_sc_hd__sdfrtp_1 c656 (.CLK(clknet_leaf_28_clk),
    .D(clknet_1_1__leaf_net530),
    .RESET_B(net320),
    .SCD(net546),
    .SCE(net550),
    .Q(net552));
 sky130_fd_sc_hd__nand3b_1 c657 (.A_N(net546),
    .B(net456),
    .C(net534),
    .Y(net553));
 sky130_fd_sc_hd__or4bb_2 c658 (.A(net740),
    .B(net221),
    .C_N(net528),
    .D_N(net699),
    .X(net554));
 sky130_fd_sc_hd__mux4_4 c659 (.A0(net553),
    .A1(net552),
    .A2(net546),
    .A3(net340),
    .S0(net529),
    .S1(net699),
    .X(net555));
 sky130_fd_sc_hd__and2b_2 c66 (.A_N(net766),
    .B(net3),
    .X(net4));
 sky130_fd_sc_hd__mux4_2 c660 (.A0(net550),
    .A1(net543),
    .A2(clknet_1_0__leaf_net547),
    .A3(net809),
    .S0(net816),
    .S1(net699),
    .X(net556));
 sky130_fd_sc_hd__nor3b_1 c661 (.A(net740),
    .B(net548),
    .C_N(net209),
    .Y(net557));
 sky130_fd_sc_hd__nor3b_1 c662 (.A(net301),
    .B(net893),
    .C_N(net413),
    .Y(net558));
 sky130_fd_sc_hd__sdfxbp_1 c663 (.CLK(clknet_leaf_31_clk),
    .D(net543),
    .SCD(net946),
    .SCE(net554),
    .Q(net559));
 sky130_fd_sc_hd__sdfsbp_1 c664 (.CLK(clknet_leaf_26_clk),
    .D(net453),
    .SCD(net871),
    .SCE(net860),
    .SET_B(net916),
    .Q(net561),
    .Q_N(net560));
 sky130_fd_sc_hd__a2111oi_1 c665 (.A1(net529),
    .A2(net552),
    .B1(net549),
    .C1(net557),
    .D1(net700),
    .Y(net562));
 sky130_fd_sc_hd__sdfsbp_1 c666 (.CLK(clknet_leaf_28_clk),
    .D(net950),
    .SCD(clknet_1_1__leaf_net530),
    .SCE(net449),
    .SET_B(net913),
    .Q(net563));
 sky130_fd_sc_hd__sdfstp_1 c667 (.CLK(clknet_leaf_31_clk),
    .D(net920),
    .SCD(net320),
    .SCE(net554),
    .SET_B(net910),
    .Q(net564));
 sky130_fd_sc_hd__or3b_1 c668 (.A(net561),
    .B(net564),
    .C_N(net548),
    .X(net565));
 sky130_fd_sc_hd__sdfstp_2 c669 (.CLK(clknet_leaf_28_clk),
    .D(net562),
    .SCD(net564),
    .SCE(net943),
    .SET_B(clknet_1_1__leaf_net670),
    .Q(net566));
 sky130_fd_sc_hd__and2_1 c67 (.A(net776),
    .B(net2),
    .X(net5));
 sky130_fd_sc_hd__nor3_1 c670 (.A(net558),
    .B(net565),
    .C(net564),
    .Y(net567));
 sky130_fd_sc_hd__or4bb_2 c671 (.A(net563),
    .B(net548),
    .C_N(net546),
    .D_N(net816),
    .X(net568));
 sky130_fd_sc_hd__sdfbbn_1 c672 (.CLK_N(clknet_leaf_28_clk),
    .D(net878),
    .RESET_B(net893),
    .SCD(clknet_1_0__leaf_net463),
    .SCE(clknet_1_1__leaf_net530),
    .SET_B(net669),
    .Q(net570),
    .Q_N(net569));
 sky130_fd_sc_hd__mux4_2 c673 (.A0(net555),
    .A1(net860),
    .A2(net450),
    .A3(net539),
    .S0(net893),
    .S1(clknet_1_1__leaf_net671),
    .X(net571));
 sky130_fd_sc_hd__sdfbbn_1 c674 (.CLK_N(clknet_leaf_28_clk),
    .D(net552),
    .RESET_B(net539),
    .SCD(clknet_1_0__leaf_net476),
    .SCE(net569),
    .SET_B(net669),
    .Q(net573),
    .Q_N(net572));
 sky130_fd_sc_hd__mux4_4 c675 (.A0(net570),
    .A1(net539),
    .A2(net893),
    .A3(net567),
    .S0(clknet_1_0__leaf_net547),
    .S1(net816),
    .X(net574));
 sky130_fd_sc_hd__sdfbbp_1 c676 (.CLK(clknet_leaf_26_clk),
    .D(net573),
    .RESET_B(net759),
    .SCD(clknet_1_0__leaf_net476),
    .SCE(net455),
    .SET_B(clknet_1_0__leaf_net672),
    .Q(net576),
    .Q_N(net575));
 sky130_fd_sc_hd__a2111oi_1 c677 (.A1(net525),
    .A2(net561),
    .B1(clknet_1_1__leaf_net547),
    .C1(net539),
    .D1(net872),
    .Y(net577));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net871),
    .A1(net569),
    .A2(net878),
    .A3(net575),
    .S0(clknet_1_0__leaf_net672),
    .S1(net702),
    .X(net578));
 sky130_fd_sc_hd__mux4_4 c679 (.A0(clknet_1_1__leaf_net463),
    .A1(net450),
    .A2(net570),
    .A3(net560),
    .S0(net525),
    .S1(net777),
    .X(net579));
 sky130_fd_sc_hd__nor2b_1 c68 (.A(net2),
    .B_N(net4),
    .Y(net6));
 sky130_fd_sc_hd__a2111o_2 c680 (.A1(net552),
    .A2(net576),
    .B1(clknet_1_1__leaf_net547),
    .C1(clknet_1_0__leaf_net577),
    .D1(net878),
    .X(net794));
 sky130_fd_sc_hd__a2111o_4 c681 (.A1(net576),
    .A2(net870),
    .B1(net872),
    .C1(clknet_1_1__leaf_net671),
    .D1(clknet_1_0__leaf_net672),
    .X(net580));
 sky130_fd_sc_hd__sdfbbn_1 c682 (.CLK_N(clknet_leaf_26_clk),
    .D(net539),
    .RESET_B(net554),
    .SCD(net573),
    .SCE(net566),
    .SET_B(net924),
    .Q(net581));
 sky130_fd_sc_hd__sdfbbn_1 c683 (.CLK_N(clknet_leaf_27_clk),
    .D(net417),
    .RESET_B(clknet_1_0__leaf_net238),
    .SCD(net860),
    .SCE(clknet_1_0__leaf_net463),
    .SET_B(net569),
    .Q(net583),
    .Q_N(net582));
 sky130_fd_sc_hd__mux4_2 c684 (.A0(net877),
    .A1(net567),
    .A2(net582),
    .A3(net860),
    .S0(clknet_1_1__leaf_net547),
    .S1(net417),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(clknet_1_1__leaf_net577),
    .A1(net580),
    .A2(net570),
    .A3(net582),
    .S0(net220),
    .S1(net575),
    .X(net585));
 sky130_fd_sc_hd__a2111o_2 c686 (.A1(net583),
    .A2(net561),
    .B1(clknet_1_0__leaf_net585),
    .C1(net573),
    .D1(net575),
    .X(net586));
 sky130_fd_sc_hd__a2111oi_1 c687 (.A1(net581),
    .A2(net784),
    .B1(net576),
    .C1(net759),
    .D1(net704),
    .Y(net587));
 sky130_fd_sc_hd__mux4_4 c688 (.A0(net587),
    .A1(clknet_1_0__leaf_net578),
    .A2(net567),
    .A3(net417),
    .S0(net449),
    .S1(clknet_1_0__leaf_net672),
    .X(net588));
 sky130_fd_sc_hd__mux4_2 c689 (.A0(clknet_1_0__leaf_net547),
    .A1(net874),
    .A2(net566),
    .A3(clknet_1_0__leaf_net794),
    .S0(net560),
    .S1(net701),
    .X(net589));
 sky130_fd_sc_hd__nor2_1 c69 (.A(net3),
    .B(net790),
    .Y(net7));
 sky130_fd_sc_hd__sdfbbp_1 c690 (.CLK(clknet_leaf_27_clk),
    .D(net583),
    .RESET_B(net860),
    .SCD(net417),
    .SCE(net945),
    .SET_B(net911),
    .Q(net590));
 sky130_fd_sc_hd__mux4_2 c691 (.A0(net589),
    .A1(net590),
    .A2(clknet_1_0__leaf_net238),
    .A3(net572),
    .S0(net784),
    .S1(net669),
    .X(net591));
 sky130_fd_sc_hd__o2111a_4 c692 (.A1(net855),
    .A2(net877),
    .B1(net314),
    .C1(net705),
    .D1(net706),
    .X(net592));
 sky130_fd_sc_hd__a2111oi_1 c693 (.A1(net564),
    .A2(net536),
    .B1(net762),
    .C1(net784),
    .D1(net896),
    .Y(net593));
 sky130_fd_sc_hd__sdfbbn_1 c694 (.CLK_N(clknet_leaf_27_clk),
    .D(clknet_1_1__leaf_net578),
    .RESET_B(clknet_1_1__leaf_net592),
    .SCD(net483),
    .SCE(clknet_1_0__leaf_net585),
    .SET_B(net863),
    .Q(net595),
    .Q_N(net594));
 sky130_fd_sc_hd__mux4_4 c695 (.A0(clknet_1_1__leaf_net585),
    .A1(net874),
    .A2(net535),
    .A3(net594),
    .S0(clknet_1_0__leaf_net142),
    .S1(net326),
    .X(net596));
 sky130_fd_sc_hd__mux4_4 c696 (.A0(net304),
    .A1(clknet_1_1__leaf_net586),
    .A2(net595),
    .A3(clknet_1_1__leaf_net585),
    .S0(net256),
    .S1(net682),
    .X(net597));
 sky130_fd_sc_hd__mux4_2 c697 (.A0(net256),
    .A1(net762),
    .A2(clknet_1_0__leaf_net476),
    .A3(net872),
    .S0(net891),
    .S1(net703),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net343),
    .A1(net593),
    .A2(net735),
    .A3(net897),
    .S0(net703),
    .S1(net704),
    .X(net599));
 sky130_fd_sc_hd__mux4_2 c699 (.A0(net595),
    .A1(net870),
    .A2(net872),
    .A3(net897),
    .S0(net891),
    .S1(net704),
    .X(net600));
 sky130_fd_sc_hd__nand2b_4 c70 (.A_N(net5),
    .B(net2),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(clknet_1_0__leaf_net597),
    .A1(net746),
    .A2(clknet_1_0__leaf_net586),
    .A3(clknet_1_0__leaf_net379),
    .S0(net343),
    .S1(net703),
    .X(net601));
 sky130_fd_sc_hd__o2111a_4 c701 (.A1(net315),
    .A2(net600),
    .B1(net566),
    .C1(clknet_1_0__leaf_net142),
    .D1(net568),
    .X(net602));
 sky130_fd_sc_hd__mux4_2 c702 (.A0(net535),
    .A1(clknet_1_0__leaf_net794),
    .A2(clknet_1_0__leaf_net476),
    .A3(net564),
    .S0(clknet_1_0__leaf_net142),
    .S1(clknet_1_1__leaf_net671),
    .X(net603));
 sky130_fd_sc_hd__sdfbbn_1 c703 (.CLK_N(clknet_leaf_23_clk),
    .D(clknet_1_0__leaf_net142),
    .RESET_B(clknet_1_1__leaf_net476),
    .SCD(net420),
    .SCE(clknet_1_1__leaf_net671),
    .SET_B(clknet_1_1__leaf_net708),
    .Q(net805),
    .Q_N(net604));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net536),
    .A1(clknet_1_1__leaf_net503),
    .A2(net220),
    .A3(net384),
    .S0(clknet_1_0__leaf_net476),
    .S1(net526),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net385),
    .A1(net256),
    .A2(net897),
    .A3(net572),
    .S0(net712),
    .S1(net714),
    .X(net606));
 sky130_fd_sc_hd__a2111oi_2 c706 (.A1(net606),
    .A2(clknet_1_0__leaf_net142),
    .B1(clknet_1_0__leaf_net708),
    .C1(net709),
    .D1(net711),
    .Y(net607));
 sky130_fd_sc_hd__mux4_2 c707 (.A0(net573),
    .A1(clknet_1_0__leaf_net503),
    .A2(net600),
    .A3(net897),
    .S0(net455),
    .S1(net710),
    .X(net608));
 sky130_fd_sc_hd__sdfbbp_1 c708 (.CLK(clknet_leaf_27_clk),
    .D(clknet_1_0__leaf_net596),
    .RESET_B(clknet_1_0__leaf_net592),
    .SCD(net874),
    .SCE(net951),
    .SET_B(net713),
    .Q(net609));
 sky130_fd_sc_hd__a2111o_1 c709 (.A1(net885),
    .A2(net607),
    .B1(net863),
    .C1(clknet_1_0__leaf_net794),
    .D1(clknet_1_1__leaf_net596),
    .X(net610));
 sky130_fd_sc_hd__or4bb_1 c71 (.A(net789),
    .B(net8),
    .C_N(net3),
    .D_N(net1),
    .X(net9));
 sky130_fd_sc_hd__mux4_2 c710 (.A0(net602),
    .A1(net885),
    .A2(net865),
    .A3(clknet_1_0__leaf_net238),
    .S0(net572),
    .S1(net682),
    .X(net611));
 sky130_fd_sc_hd__mux4_4 c711 (.A0(net526),
    .A1(net600),
    .A2(clknet_1_0__leaf_net142),
    .A3(net566),
    .S0(clknet_1_1__leaf_net597),
    .S1(net710),
    .X(net612));
 sky130_fd_sc_hd__mux4_4 c712 (.A0(net566),
    .A1(clknet_1_1__leaf_net610),
    .A2(net784),
    .A3(net220),
    .S0(net700),
    .S1(net715),
    .X(net613));
 sky130_fd_sc_hd__sdfbbn_1 c713 (.CLK_N(clknet_leaf_23_clk),
    .D(clknet_1_0__leaf_net794),
    .RESET_B(clknet_1_0__leaf_net610),
    .SCD(net930),
    .SCE(net714),
    .SET_B(net718),
    .Q(net614));
 sky130_fd_sc_hd__mux4_2 c714 (.A0(net881),
    .A1(clknet_1_0__leaf_net289),
    .A2(net865),
    .A3(net456),
    .S0(net732),
    .S1(clknet_1_0__leaf_net707),
    .X(net615));
 sky130_fd_sc_hd__mux4_2 c715 (.A0(clknet_1_0__leaf_net238),
    .A1(clknet_1_1__leaf_net615),
    .A2(net483),
    .A3(net746),
    .S0(net455),
    .S1(net698),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net508),
    .A1(net398),
    .A2(clknet_1_0__leaf_net238),
    .A3(clknet_1_0__leaf_net615),
    .S0(net816),
    .S1(net719),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net456),
    .A1(net496),
    .A2(net897),
    .A3(net826),
    .S0(net865),
    .S1(net716),
    .X(net618));
 sky130_fd_sc_hd__mux4_2 c718 (.A0(net609),
    .A1(net864),
    .A2(net496),
    .A3(net809),
    .S0(clknet_1_0__leaf_net691),
    .S1(net700),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net221),
    .A1(net870),
    .A2(net604),
    .A3(net511),
    .S0(net698),
    .S1(net720),
    .X(net620));
 sky130_fd_sc_hd__nand2b_2 c72 (.A_N(net9),
    .B(net4),
    .Y(net10));
 sky130_fd_sc_hd__mux4_2 c720 (.A0(net511),
    .A1(clknet_1_0__leaf_net615),
    .A2(clknet_1_0__leaf_net619),
    .A3(net874),
    .S0(net865),
    .S1(net891),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net496),
    .A1(net398),
    .A2(clknet_1_1__leaf_net794),
    .A3(net697),
    .S0(net700),
    .S1(net719),
    .X(net622));
 sky130_fd_sc_hd__mux4_4 c722 (.A0(net614),
    .A1(clknet_1_0__leaf_net610),
    .A2(net874),
    .A3(clknet_1_0__leaf_net379),
    .S0(net826),
    .S1(net893),
    .X(net623));
 sky130_fd_sc_hd__mux4_2 c723 (.A0(clknet_1_0__leaf_net513),
    .A1(clknet_1_0__leaf_net489),
    .A2(clknet_1_1__leaf_net794),
    .A3(net881),
    .S0(clknet_1_0__leaf_net691),
    .S1(clknet_1_0__leaf_net707),
    .X(net624));
 sky130_fd_sc_hd__mux4_2 c724 (.A0(net483),
    .A1(clknet_1_0__leaf_net513),
    .A2(clknet_1_1__leaf_net489),
    .A3(net863),
    .S0(clknet_1_1__leaf_net794),
    .S1(clknet_1_1__leaf_net691),
    .X(net625));
 sky130_fd_sc_hd__mux4_2 c725 (.A0(net568),
    .A1(net622),
    .A2(clknet_1_0__leaf_net379),
    .A3(net385),
    .S0(net420),
    .S1(net456),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net864),
    .A1(clknet_1_1__leaf_net476),
    .A2(net870),
    .A3(net881),
    .S0(net722),
    .S1(net723),
    .X(net627));
 sky130_fd_sc_hd__mux4_2 c727 (.A0(net326),
    .A1(clknet_1_1__leaf_net794),
    .A2(net784),
    .A3(net698),
    .S0(net717),
    .S1(net721),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net620),
    .A1(clknet_1_1__leaf_net794),
    .A2(net865),
    .A3(net398),
    .S0(net723),
    .S1(net724),
    .X(net629));
 sky130_fd_sc_hd__mux4_2 c729 (.A0(clknet_1_0__leaf_net379),
    .A1(clknet_1_1__leaf_net619),
    .A2(net398),
    .A3(clknet_1_0__leaf_net289),
    .S0(clknet_1_0__leaf_net238),
    .S1(net725),
    .X(net630));
 sky130_fd_sc_hd__nor2_2 c73 (.A(net5),
    .B(net772),
    .Y(net11));
 sky130_fd_sc_hd__mux4_2 c730 (.A0(net746),
    .A1(net511),
    .A2(clknet_1_1__leaf_net707),
    .A3(clknet_1_1__leaf_net726),
    .S0(net727),
    .S1(net728),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(clknet_1_1__leaf_net476),
    .A1(clknet_1_0__leaf_net631),
    .A2(net784),
    .A3(net722),
    .S0(net723),
    .S1(clknet_1_0__leaf_net726),
    .X(net632));
 sky130_fd_sc_hd__mux4_2 c732 (.A0(clknet_1_1__leaf_net631),
    .A1(clknet_1_1__leaf_net794),
    .A2(clknet_1_0__leaf_net238),
    .A3(net719),
    .S0(clknet_1_0__leaf_net726),
    .S1(net729),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net886),
    .A1(net618),
    .A2(net628),
    .A3(clknet_1_1__leaf_net794),
    .S0(net865),
    .S1(clknet_1_0__leaf_net631),
    .X(net634));
 sky130_fd_sc_hd__mux4_4 c734 (.A0(clknet_1_1__leaf_net489),
    .A1(net456),
    .A2(clknet_1_1__leaf_net631),
    .A3(net326),
    .S0(net730),
    .S1(net731),
    .X(net635));
 sky130_fd_sc_hd__nor2_1 c74 (.A(net1),
    .B(net9),
    .Y(net12));
 sky130_fd_sc_hd__nand2_8 c75 (.A(net4),
    .B(net3),
    .Y(net13));
 sky130_fd_sc_hd__or2_4 c76 (.A(net763),
    .B(net0),
    .X(net14));
 sky130_fd_sc_hd__and2_4 c77 (.A(net13),
    .B(net751),
    .X(net15));
 sky130_fd_sc_hd__o2111ai_4 c78 (.A1(net11),
    .A2(net758),
    .B1(net767),
    .C1(net13),
    .D1(net15),
    .Y(net16));
 sky130_fd_sc_hd__nand2_1 c79 (.A(net8),
    .B(net14),
    .Y(net17));
 sky130_fd_sc_hd__and2_4 c80 (.A(net16),
    .B(net732),
    .X(net18));
 sky130_fd_sc_hd__o2111ai_4 c81 (.A1(net772),
    .A2(net7),
    .B1(net18),
    .C1(net15),
    .D1(net14),
    .Y(net19));
 sky130_fd_sc_hd__or4bb_4 c82 (.A(net17),
    .B(net15),
    .C_N(net5),
    .D_N(net14),
    .X(net20));
 sky130_fd_sc_hd__mux4_2 c83 (.A0(net16),
    .A1(net17),
    .A2(net20),
    .A3(net14),
    .S0(net13),
    .S1(net19),
    .X(net21));
 sky130_fd_sc_hd__or2b_1 c84 (.A(net16),
    .B_N(net14),
    .X(net22));
 sky130_fd_sc_hd__and2b_1 c85 (.A_N(net2),
    .B(net4),
    .X(net23));
 sky130_fd_sc_hd__or2_1 c86 (.A(net780),
    .B(net16),
    .X(net24));
 sky130_fd_sc_hd__nand2b_4 c87 (.A_N(net750),
    .B(net735),
    .Y(net25));
 sky130_fd_sc_hd__or4bb_1 c88 (.A(net24),
    .B(net14),
    .C_N(net12),
    .D_N(net8),
    .X(net26));
 sky130_fd_sc_hd__and2_0 c89 (.A(net4),
    .B(net25),
    .X(net27));
 sky130_fd_sc_hd__and2_1 c90 (.A(net6),
    .B(net25),
    .X(net28));
 sky130_fd_sc_hd__nand2_1 c91 (.A(net781),
    .B(net23),
    .Y(net29));
 sky130_fd_sc_hd__or2_1 c92 (.A(net758),
    .B(net778),
    .X(net30));
 sky130_fd_sc_hd__or2_2 c93 (.A(net22),
    .B(net25),
    .X(net31));
 sky130_fd_sc_hd__nand2_1 c94 (.A(net25),
    .B(net28),
    .Y(net32));
 sky130_fd_sc_hd__and2_2 c95 (.A(net29),
    .B(net25),
    .X(net33));
 sky130_fd_sc_hd__o2111a_2 c96 (.A1(net27),
    .A2(net33),
    .B1(net4),
    .C1(net746),
    .D1(net28),
    .X(net34));
 sky130_fd_sc_hd__mux4_2 c97 (.A0(net31),
    .A1(net13),
    .A2(net6),
    .A3(net24),
    .S0(net25),
    .S1(net30),
    .X(net839));
 sky130_fd_sc_hd__or2b_1 c98 (.A(net7),
    .B_N(net31),
    .X(net35));
 sky130_fd_sc_hd__nor2_2 c99 (.A(net28),
    .B(net33),
    .Y(net36));
 sky130_fd_sc_hd__sdfstp_1 merge740 (.CLK(clknet_leaf_32_clk),
    .D(net199),
    .SCD(net320),
    .SCE(net197),
    .SET_B(net316),
    .Q(net636));
 sky130_fd_sc_hd__dfxbp_1 s741 (.CLK(clknet_leaf_13_clk),
    .D(net56),
    .Q(net847),
    .Q_N(net637));
 sky130_fd_sc_hd__dfxbp_1 s742 (.CLK(clknet_leaf_13_clk),
    .D(net60),
    .Q(net824),
    .Q_N(net638));
 sky130_fd_sc_hd__dfxtp_1 s743 (.CLK(clknet_leaf_6_clk),
    .D(net103),
    .Q(net639));
 sky130_fd_sc_hd__dfxtp_1 s744 (.CLK(clknet_leaf_6_clk),
    .D(net105),
    .Q(net640));
 sky130_fd_sc_hd__dfxtp_1 s745 (.CLK(clknet_leaf_7_clk),
    .D(net126),
    .Q(net641));
 sky130_fd_sc_hd__dlclkp_1 s746 (.CLK(clknet_leaf_7_clk),
    .GATE(net129),
    .GCLK(net642));
 sky130_fd_sc_hd__dlclkp_2 s747 (.CLK(clknet_leaf_7_clk),
    .GATE(net131),
    .GCLK(net643));
 sky130_fd_sc_hd__dlclkp_4 s748 (.CLK(clknet_leaf_14_clk),
    .GATE(net177),
    .GCLK(net798));
 sky130_fd_sc_hd__dlxbn_1 s749 (.D(net216),
    .GATE_N(clknet_leaf_3_clk),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__dlxbn_2 s750 (.D(net223),
    .GATE_N(clknet_leaf_8_clk),
    .Q(net809),
    .Q_N(net646));
 sky130_fd_sc_hd__dlxbp_1 s751 (.D(net224),
    .GATE(clknet_leaf_8_clk),
    .Q(net648),
    .Q_N(net647));
 sky130_fd_sc_hd__dlxtn_1 s752 (.D(net242),
    .GATE_N(clknet_leaf_7_clk),
    .Q(net803));
 sky130_fd_sc_hd__dlxtn_1 s753 (.D(net243),
    .GATE_N(clknet_leaf_8_clk),
    .Q(net649));
 sky130_fd_sc_hd__dlxtn_1 s754 (.D(net263),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net650));
 sky130_fd_sc_hd__dlxtp_1 s755 (.D(net272),
    .GATE(clknet_leaf_10_clk),
    .Q(net800));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s756 (.D(net273),
    .SLEEP_B(clknet_leaf_18_clk),
    .Q(net651));
 sky130_fd_sc_hd__dfxbp_1 s757 (.CLK(clknet_leaf_18_clk),
    .D(net292),
    .Q(net822),
    .Q_N(net652));
 sky130_fd_sc_hd__dfxbp_1 s758 (.CLK(clknet_leaf_15_clk),
    .D(net293),
    .Q(net838),
    .Q_N(net653));
 sky130_fd_sc_hd__dfxtp_1 s759 (.CLK(clknet_leaf_15_clk),
    .D(net294),
    .Q(net851));
 sky130_fd_sc_hd__dfxtp_1 s760 (.CLK(clknet_leaf_15_clk),
    .D(net295),
    .Q(net836));
 sky130_fd_sc_hd__dfxtp_1 s761 (.CLK(clknet_leaf_16_clk),
    .D(net296),
    .Q(net846));
 sky130_fd_sc_hd__dlclkp_1 s762 (.CLK(clknet_leaf_16_clk),
    .GATE(net297),
    .GCLK(net841));
 sky130_fd_sc_hd__dlclkp_2 s763 (.CLK(clknet_leaf_32_clk),
    .GATE(net368),
    .GCLK(net814));
 sky130_fd_sc_hd__dlclkp_4 s764 (.CLK(clknet_leaf_19_clk),
    .GATE(net382),
    .GCLK(net654));
 sky130_fd_sc_hd__dlxbn_1 s765 (.D(net383),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net656),
    .Q_N(net655));
 sky130_fd_sc_hd__dlxbn_1 s766 (.D(net386),
    .GATE_N(clknet_leaf_17_clk),
    .Q(net658),
    .Q_N(net657));
 sky130_fd_sc_hd__dlxbp_1 s767 (.D(net387),
    .GATE(clknet_leaf_19_clk),
    .Q(net660),
    .Q_N(net659));
 sky130_fd_sc_hd__dlxtn_1 s768 (.D(net389),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net661));
 sky130_fd_sc_hd__dlxtn_1 s769 (.D(net390),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net662));
 sky130_fd_sc_hd__dlxtn_1 s770 (.D(net391),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net663));
 sky130_fd_sc_hd__dlxtp_1 s771 (.D(net392),
    .GATE(clknet_leaf_20_clk),
    .Q(net664));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s772 (.D(net400),
    .SLEEP_B(clknet_leaf_17_clk),
    .Q(net665));
 sky130_fd_sc_hd__dfxbp_1 s773 (.CLK(clknet_leaf_20_clk),
    .D(net402),
    .Q(net802),
    .Q_N(net666));
 sky130_fd_sc_hd__dfxbp_1 s774 (.CLK(clknet_leaf_17_clk),
    .D(net403),
    .Q(net667));
 sky130_fd_sc_hd__dfxtp_1 s775 (.CLK(clknet_leaf_17_clk),
    .D(net404),
    .Q(net828));
 sky130_fd_sc_hd__dfxtp_1 s776 (.CLK(clknet_leaf_17_clk),
    .D(net405),
    .Q(net668));
 sky130_fd_sc_hd__dfxtp_2 s777 (.CLK(clknet_leaf_32_clk),
    .D(net427),
    .Q(net669));
 sky130_fd_sc_hd__dlclkp_1 s778 (.CLK(clknet_leaf_31_clk),
    .GATE(net431),
    .GCLK(net670));
 sky130_fd_sc_hd__dlclkp_2 s779 (.CLK(clknet_leaf_1_clk),
    .GATE(net464),
    .GCLK(net671));
 sky130_fd_sc_hd__dlclkp_4 s780 (.CLK(clknet_leaf_25_clk),
    .GATE(net473),
    .GCLK(net672));
 sky130_fd_sc_hd__dlxbn_1 s781 (.D(net475),
    .GATE_N(clknet_leaf_1_clk),
    .Q(net673));
 sky130_fd_sc_hd__dlxbn_1 s782 (.D(net477),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__dlxbp_1 s783 (.D(net478),
    .GATE(clknet_leaf_25_clk),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dlxtn_1 s784 (.D(net480),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net678));
 sky130_fd_sc_hd__dlxtn_1 s785 (.D(net481),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net679));
 sky130_fd_sc_hd__dlxtn_1 s786 (.D(net488),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net680));
 sky130_fd_sc_hd__dlxtp_1 s787 (.D(net495),
    .GATE(clknet_leaf_19_clk),
    .Q(net681));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s788 (.D(net497),
    .SLEEP_B(clknet_leaf_24_clk),
    .Q(net682));
 sky130_fd_sc_hd__dfxbp_1 s789 (.CLK(clknet_leaf_24_clk),
    .D(net499),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__dfxbp_1 s790 (.CLK(clknet_leaf_19_clk),
    .D(net500),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__dfxtp_1 s791 (.CLK(clknet_leaf_24_clk),
    .D(net502),
    .Q(net687));
 sky130_fd_sc_hd__dfxtp_2 s792 (.CLK(clknet_leaf_20_clk),
    .D(net507),
    .Q(net688));
 sky130_fd_sc_hd__dfxtp_1 s793 (.CLK(clknet_leaf_21_clk),
    .D(net509),
    .Q(net806));
 sky130_fd_sc_hd__dlclkp_1 s794 (.CLK(clknet_leaf_20_clk),
    .GATE(net510),
    .GCLK(net689));
 sky130_fd_sc_hd__dlclkp_2 s795 (.CLK(clknet_leaf_20_clk),
    .GATE(net515),
    .GCLK(net690));
 sky130_fd_sc_hd__dlclkp_4 s796 (.CLK(clknet_leaf_20_clk),
    .GATE(net516),
    .GCLK(net691));
 sky130_fd_sc_hd__dlxbn_1 s797 (.D(net518),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net693),
    .Q_N(net692));
 sky130_fd_sc_hd__dlxbn_1 s798 (.D(net519),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net797),
    .Q_N(net694));
 sky130_fd_sc_hd__dlxbp_1 s799 (.D(net520),
    .GATE(clknet_leaf_20_clk),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__dlxtn_1 s800 (.D(net521),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net697));
 sky130_fd_sc_hd__dlxtn_1 s801 (.D(net523),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net698));
 sky130_fd_sc_hd__dlxtn_2 s802 (.D(net544),
    .GATE_N(clknet_leaf_29_clk),
    .Q(net816));
 sky130_fd_sc_hd__dlxtp_1 s803 (.D(net545),
    .GATE(clknet_leaf_28_clk),
    .Q(net699));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s804 (.D(net556),
    .SLEEP_B(clknet_leaf_28_clk),
    .Q(net700));
 sky130_fd_sc_hd__dfxbp_1 s805 (.CLK(clknet_leaf_27_clk),
    .D(net571),
    .Q(net701));
 sky130_fd_sc_hd__dfxbp_1 s806 (.CLK(clknet_leaf_27_clk),
    .D(net574),
    .Q(net702));
 sky130_fd_sc_hd__dfxtp_1 s807 (.CLK(clknet_leaf_26_clk),
    .D(net579),
    .Q(net703));
 sky130_fd_sc_hd__dfxtp_1 s808 (.CLK(clknet_leaf_27_clk),
    .D(net584),
    .Q(net704));
 sky130_fd_sc_hd__dfxtp_1 s809 (.CLK(clknet_leaf_27_clk),
    .D(net588),
    .Q(net705));
 sky130_fd_sc_hd__dlclkp_1 s810 (.CLK(clknet_leaf_27_clk),
    .GATE(net591),
    .GCLK(net706));
 sky130_fd_sc_hd__dlclkp_2 s811 (.CLK(clknet_leaf_25_clk),
    .GATE(net598),
    .GCLK(net707));
 sky130_fd_sc_hd__dlclkp_4 s812 (.CLK(clknet_leaf_23_clk),
    .GATE(net599),
    .GCLK(net708));
 sky130_fd_sc_hd__dlxbn_1 s813 (.D(net601),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net710),
    .Q_N(net709));
 sky130_fd_sc_hd__dlxbn_1 s814 (.D(net603),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__dlxbp_1 s815 (.D(net605),
    .GATE(clknet_leaf_23_clk),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__dlxtn_1 s816 (.D(net608),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net715));
 sky130_fd_sc_hd__dlxtn_1 s817 (.D(net611),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net716));
 sky130_fd_sc_hd__dlxtn_1 s818 (.D(net612),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net717));
 sky130_fd_sc_hd__dlxtp_1 s819 (.D(net613),
    .GATE(clknet_leaf_23_clk),
    .Q(net718));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s820 (.D(net616),
    .SLEEP_B(clknet_leaf_24_clk),
    .Q(net719));
 sky130_fd_sc_hd__dfxbp_1 s821 (.CLK(clknet_leaf_24_clk),
    .D(net617),
    .Q(net720));
 sky130_fd_sc_hd__dfxbp_1 s822 (.CLK(clknet_leaf_22_clk),
    .D(net621),
    .Q(net721));
 sky130_fd_sc_hd__dfxtp_1 s823 (.CLK(clknet_leaf_23_clk),
    .D(net623),
    .Q(net722));
 sky130_fd_sc_hd__dfxtp_1 s824 (.CLK(clknet_leaf_22_clk),
    .D(net624),
    .Q(net723));
 sky130_fd_sc_hd__dfxtp_1 s825 (.CLK(clknet_leaf_22_clk),
    .D(net625),
    .Q(net724));
 sky130_fd_sc_hd__dlclkp_1 s826 (.CLK(clknet_leaf_24_clk),
    .GATE(net626),
    .GCLK(net725));
 sky130_fd_sc_hd__dlclkp_2 s827 (.CLK(clknet_leaf_22_clk),
    .GATE(net627),
    .GCLK(net726));
 sky130_fd_sc_hd__dlclkp_4 s828 (.CLK(clknet_leaf_21_clk),
    .GATE(net629),
    .GCLK(net727));
 sky130_fd_sc_hd__dlxbn_1 s829 (.D(net630),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net728));
 sky130_fd_sc_hd__dlxbn_1 s830 (.D(net632),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net729));
 sky130_fd_sc_hd__dlxbp_1 s831 (.D(net633),
    .GATE(clknet_leaf_22_clk),
    .Q(net730));
 sky130_fd_sc_hd__dlxtn_1 s832 (.D(net634),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net731));
 sky130_fd_sc_hd__dlxtn_2 s833 (.D(net635),
    .GATE_N(clknet_leaf_22_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(in0),
    .X(net732));
 sky130_fd_sc_hd__buf_4 input2 (.A(in1),
    .X(net733));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(in11),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net736));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(in13),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net738));
 sky130_fd_sc_hd__buf_2 input8 (.A(in15),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in16),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net742));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net743));
 sky130_fd_sc_hd__buf_1 input13 (.A(in2),
    .X(net744));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net746));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(in22),
    .X(net747));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net749));
 sky130_fd_sc_hd__buf_2 input19 (.A(in25),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in26),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(in27),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net753));
 sky130_fd_sc_hd__buf_1 input23 (.A(net912),
    .X(net754));
 sky130_fd_sc_hd__buf_6 input24 (.A(in3),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(in31),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net758));
 sky130_fd_sc_hd__buf_4 input28 (.A(in33),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(in35),
    .X(net761));
 sky130_fd_sc_hd__buf_2 input31 (.A(in36),
    .X(net762));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(in38),
    .X(net764));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(in39),
    .X(net765));
 sky130_fd_sc_hd__buf_2 input35 (.A(in4),
    .X(net766));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net767));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(in42),
    .X(net769));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(in44),
    .X(net771));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(in45),
    .X(net772));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(in47),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(in48),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in49),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(in5),
    .X(net777));
 sky130_fd_sc_hd__buf_2 input47 (.A(in50),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(in52),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net781));
 sky130_fd_sc_hd__buf_6 input51 (.A(in54),
    .X(net782));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(in55),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_8 input53 (.A(in56),
    .X(net784));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(in58),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(in59),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(in6),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(in60),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(in61),
    .X(net790));
 sky130_fd_sc_hd__buf_12 input60 (.A(in7),
    .X(net791));
 sky130_fd_sc_hd__buf_1 input61 (.A(in8),
    .X(net792));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(in9),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(clknet_1_0__leaf_net794),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output64 (.A(net795),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(clknet_1_1__leaf_net796),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net797),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net798),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output68 (.A(net799),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net800),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(clknet_1_1__leaf_net801),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net802),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net803),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net804),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output74 (.A(net805),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output75 (.A(net806),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output76 (.A(net807),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net808),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output78 (.A(net809),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output79 (.A(net810),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output80 (.A(net811),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(clknet_1_1__leaf_net812),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output82 (.A(net813),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net814),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(clknet_1_1__leaf_net815),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output85 (.A(net816),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net817),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_1__leaf_net818),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net819),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output89 (.A(net820),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output90 (.A(net821),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output91 (.A(net822),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(clknet_1_1__leaf_net823),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net824),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output94 (.A(net825),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output95 (.A(net860),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output96 (.A(net827),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output97 (.A(net828),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(clknet_1_1__leaf_net829),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output99 (.A(net830),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output100 (.A(net831),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output101 (.A(net832),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output102 (.A(net833),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(clknet_1_0__leaf_net834),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(clknet_1_1__leaf_net835),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output105 (.A(net836),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output106 (.A(net874),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output107 (.A(net838),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net839),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output109 (.A(net840),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net841),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net842),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(clknet_1_0__leaf_net843),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net844),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output114 (.A(net845),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output115 (.A(net846),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net847),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(clknet_1_1__leaf_net848),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net849),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net850),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output120 (.A(net851),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(clknet_1_1__leaf_net852),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_2 max_cap122 (.A(net465),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_1 max_cap123 (.A(net955),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_2 max_cap124 (.A(net527),
    .X(net855));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire125 (.A(net857),
    .X(net856));
 sky130_fd_sc_hd__buf_1 max_cap126 (.A(net858),
    .X(net857));
 sky130_fd_sc_hd__buf_1 max_cap127 (.A(net799),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_1 max_cap128 (.A(net421),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net826),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net863),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net863),
    .X(net862));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net326),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_2 max_cap133 (.A(net276),
    .X(net864));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net795),
    .X(net865));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap135 (.A(net96),
    .X(net866));
 sky130_fd_sc_hd__buf_1 max_cap136 (.A(net313),
    .X(net867));
 sky130_fd_sc_hd__buf_2 max_cap137 (.A(net310),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_1 max_cap138 (.A(net312),
    .X(net869));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net85),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_1 max_cap140 (.A(net557),
    .X(net871));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net873),
    .X(net872));
 sky130_fd_sc_hd__buf_6 fanout142 (.A(net874),
    .X(net873));
 sky130_fd_sc_hd__buf_6 fanout143 (.A(net837),
    .X(net874));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire144 (.A(net957),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_1 max_cap145 (.A(net958),
    .X(net876));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net191),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net112),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_2 wire148 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap149 (.A(net81),
    .X(net880));
 sky130_fd_sc_hd__buf_2 fanout150 (.A(net34),
    .X(net881));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(net84),
    .X(net882));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net188),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_2 max_cap153 (.A(net72),
    .X(net884));
 sky130_fd_sc_hd__buf_1 wire154 (.A(net959),
    .X(net885));
 sky130_fd_sc_hd__buf_4 fanout155 (.A(net370),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_1 max_cap156 (.A(net960),
    .X(net887));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire157 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire158 (.A(net890),
    .X(net889));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire159 (.A(net962),
    .X(net890));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(net800),
    .X(net891));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(net803),
    .X(net892));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net420),
    .X(net893));
 sky130_fd_sc_hd__buf_1 max_cap163 (.A(net65),
    .X(net894));
 sky130_fd_sc_hd__buf_8 fanout164 (.A(net896),
    .X(net895));
 sky130_fd_sc_hd__buf_12 fanout165 (.A(net898),
    .X(net896));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(net898),
    .X(net897));
 sky130_fd_sc_hd__buf_6 fanout167 (.A(net741),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net631 (.A(net631),
    .X(clknet_0_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net631 (.A(clknet_0_net631),
    .X(clknet_1_0__leaf_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net631 (.A(clknet_0_net631),
    .X(clknet_1_1__leaf_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net726 (.A(net726),
    .X(clknet_0_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_0__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_1__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net708 (.A(net708),
    .X(clknet_0_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_0__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_1__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net610 (.A(net610),
    .X(clknet_0_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_0__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_1__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net707 (.A(net707),
    .X(clknet_0_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_0__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_1__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net615 (.A(net615),
    .X(clknet_0_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net592 (.A(net592),
    .X(clknet_0_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_0__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_1__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net691 (.A(net691),
    .X(clknet_0_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net691 (.A(clknet_0_net691),
    .X(clknet_1_0__leaf_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net691 (.A(clknet_0_net691),
    .X(clknet_1_1__leaf_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net619 (.A(net619),
    .X(clknet_0_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net619 (.A(clknet_0_net619),
    .X(clknet_1_0__leaf_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net619 (.A(clknet_0_net619),
    .X(clknet_1_1__leaf_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net690 (.A(net690),
    .X(clknet_0_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net690 (.A(clknet_0_net690),
    .X(clknet_1_0__leaf_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net690 (.A(clknet_0_net690),
    .X(clknet_1_1__leaf_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net689 (.A(net689),
    .X(clknet_0_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net513 (.A(net513),
    .X(clknet_0_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_0__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_1__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net672 (.A(net672),
    .X(clknet_0_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net585 (.A(net585),
    .X(clknet_0_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_0__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_1__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net597 (.A(net597),
    .X(clknet_0_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_0__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_1__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net586 (.A(net586),
    .X(clknet_0_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_0__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_1__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net578 (.A(net578),
    .X(clknet_0_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net578 (.A(clknet_0_net578),
    .X(clknet_1_0__leaf_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net578 (.A(clknet_0_net578),
    .X(clknet_1_1__leaf_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net476 (.A(net476),
    .X(clknet_0_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net474 (.A(net474),
    .X(clknet_0_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_0__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_1__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net671 (.A(net671),
    .X(clknet_0_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net670 (.A(net670),
    .X(clknet_0_net670));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net670 (.A(clknet_0_net670),
    .X(clknet_1_0__leaf_net670));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net670 (.A(clknet_0_net670),
    .X(clknet_1_1__leaf_net670));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net547 (.A(net547),
    .X(clknet_0_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net794 (.A(net794),
    .X(clknet_0_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net530 (.A(net530),
    .X(clknet_0_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_0__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_1__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net439 (.A(net439),
    .X(clknet_0_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_0__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_1__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net643 (.A(net643),
    .X(clknet_0_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_0__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_1__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net228 (.A(net228),
    .X(clknet_0_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_0__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_1__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net238 (.A(net238),
    .X(clknet_0_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net235 (.A(net235),
    .X(clknet_0_net235));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net235 (.A(clknet_0_net235),
    .X(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net235 (.A(clknet_0_net235),
    .X(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net241 (.A(net241),
    .X(clknet_0_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_1__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net240 (.A(net240),
    .X(clknet_0_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net240 (.A(clknet_0_net240),
    .X(clknet_1_0__leaf_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net240 (.A(clknet_0_net240),
    .X(clknet_1_1__leaf_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net237 (.A(net237),
    .X(clknet_0_net237));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net237 (.A(clknet_0_net237),
    .X(clknet_1_0__leaf_net237));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net237 (.A(clknet_0_net237),
    .X(clknet_1_1__leaf_net237));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net249 (.A(net249),
    .X(clknet_0_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_0__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_1__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net250 (.A(net250),
    .X(clknet_0_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_0__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_1__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net236 (.A(net236),
    .X(clknet_0_net236));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net236 (.A(clknet_0_net236),
    .X(clknet_1_0__leaf_net236));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net236 (.A(clknet_0_net236),
    .X(clknet_1_1__leaf_net236));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net642 (.A(net642),
    .X(clknet_0_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net642 (.A(clknet_0_net642),
    .X(clknet_1_0__leaf_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net642 (.A(clknet_0_net642),
    .X(clknet_1_1__leaf_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net143 (.A(net143),
    .X(clknet_0_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_0__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_1__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net146 (.A(net146),
    .X(clknet_0_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net146 (.A(clknet_0_net146),
    .X(clknet_1_0__leaf_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net146 (.A(clknet_0_net146),
    .X(clknet_1_1__leaf_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net815 (.A(net815),
    .X(clknet_0_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net815 (.A(clknet_0_net815),
    .X(clknet_1_0__leaf_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net815 (.A(clknet_0_net815),
    .X(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net514 (.A(net514),
    .X(clknet_0_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net514 (.A(clknet_0_net514),
    .X(clknet_1_0__leaf_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net514 (.A(clknet_0_net514),
    .X(clknet_1_1__leaf_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net835 (.A(net835),
    .X(clknet_0_net835));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net835 (.A(clknet_0_net835),
    .X(clknet_1_0__leaf_net835));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net835 (.A(clknet_0_net835),
    .X(clknet_1_1__leaf_net835));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net834 (.A(net834),
    .X(clknet_0_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_0__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net145 (.A(net145),
    .X(clknet_0_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_1__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net286 (.A(net286),
    .X(clknet_0_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_0__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_1__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net165 (.A(net165),
    .X(clknet_0_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net166 (.A(net166),
    .X(clknet_0_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_1__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net796 (.A(net796),
    .X(clknet_0_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_0__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_1__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net829 (.A(net829),
    .X(clknet_0_net829));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net829 (.A(clknet_0_net829),
    .X(clknet_1_0__leaf_net829));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net829 (.A(clknet_0_net829),
    .X(clknet_1_1__leaf_net829));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net852 (.A(net852),
    .X(clknet_0_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net852 (.A(clknet_0_net852),
    .X(clknet_1_0__leaf_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net852 (.A(clknet_0_net852),
    .X(clknet_1_1__leaf_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net394 (.A(net394),
    .X(clknet_0_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_0__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_1__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net169 (.A(net169),
    .X(clknet_0_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net150 (.A(net150),
    .X(clknet_0_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net150 (.A(clknet_0_net150),
    .X(clknet_1_0__leaf_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net150 (.A(clknet_0_net150),
    .X(clknet_1_1__leaf_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net843 (.A(net843),
    .X(clknet_0_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net378 (.A(net378),
    .X(clknet_0_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_1__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net381 (.A(net381),
    .X(clknet_0_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_0__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_1__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net379 (.A(net379),
    .X(clknet_0_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_1__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net148 (.A(net148),
    .X(clknet_0_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net148 (.A(clknet_0_net148),
    .X(clknet_1_0__leaf_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net148 (.A(clknet_0_net148),
    .X(clknet_1_1__leaf_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net155 (.A(net155),
    .X(clknet_0_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net155 (.A(net908),
    .X(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net164 (.A(net164),
    .X(clknet_0_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_1__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net812 (.A(net812),
    .X(clknet_0_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net812 (.A(clknet_0_net812),
    .X(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net812 (.A(clknet_0_net812),
    .X(clknet_1_1__leaf_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net503 (.A(net503),
    .X(clknet_0_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_1__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net501 (.A(net501),
    .X(clknet_0_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_0__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_1__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net491 (.A(net491),
    .X(clknet_0_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_0__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net823 (.A(net823),
    .X(clknet_0_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net261 (.A(net261),
    .X(clknet_0_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net260 (.A(net260),
    .X(clknet_0_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_0__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_1__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net149 (.A(net149),
    .X(clknet_0_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net149 (.A(clknet_0_net149),
    .X(clknet_1_0__leaf_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net149 (.A(clknet_0_net149),
    .X(clknet_1_1__leaf_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net147 (.A(net147),
    .X(clknet_0_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net170 (.A(net170),
    .X(clknet_0_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_0__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_1__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net848 (.A(net848),
    .X(clknet_0_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net848 (.A(clknet_0_net848),
    .X(clknet_1_0__leaf_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net848 (.A(clknet_0_net848),
    .X(clknet_1_1__leaf_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net818 (.A(net818),
    .X(clknet_0_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net818 (.A(clknet_0_net818),
    .X(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net818 (.A(clknet_0_net818),
    .X(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net801 (.A(net801),
    .X(clknet_0_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net801 (.A(clknet_0_net801),
    .X(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net801 (.A(clknet_0_net801),
    .X(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net144 (.A(net144),
    .X(clknet_0_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_0__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_1__leaf_net144));
 sky130_fd_sc_hd__and3b_1 clone1 (.A_N(net755),
    .B(net19),
    .C(net10),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net76),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net900),
    .X(net901));
 sky130_fd_sc_hd__nand2b_1 clone4 (.A_N(net791),
    .B(net733),
    .Y(net902));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net898),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net903),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_1 clone7 (.A(clknet_0_net142),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__and3_1 clone9 (.A(net970),
    .B(net742),
    .C(net734),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(clknet_0_net155),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(clknet_1_0__leaf_net155),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net340),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net705),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(in29),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net699),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net319),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net639),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net700),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net315),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net314),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net346),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net559),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net281),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net636),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net118),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net646),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net268),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net444),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net337),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net257),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net357),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net712),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net659),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net252),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net461),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net62),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net178),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net437),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net123),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net215),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net355),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net124),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net345),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net285),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net546),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net466),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net703),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net301),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net438),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net333),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net436),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net551),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net704),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net669),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net318),
    .X(net953));
 sky130_fd_sc_hd__buf_1 max_cap1 (.A(net465),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_1 wire2 (.A(net331),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_1 wire3 (.A(net329),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_1 wire4 (.A(net222),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_1 max_cap5 (.A(net193),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_1 max_cap6 (.A(net593),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_1 max_cap7 (.A(net134),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_1 max_cap8 (.A(net962),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_1 wire9 (.A(net71),
    .X(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold14_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_D_N (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_Y (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_DE (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_D (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_SCE (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_SCD (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_D (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_SET_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_RESET_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A3 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_Q_N (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_RESET_B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_Q (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_S0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_C1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_Y (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_D1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A3 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_Y (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_B_N (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A3 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_D_N (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_D1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_D1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_X (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_SCD (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_C_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_C (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_B_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_X (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_D1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SCE (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_Y (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A3 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_S1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_RESET_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_DE (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SET_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_C (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_C (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_C (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Q_N (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A_N (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_C_N (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Q (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_C_N (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_D (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_C_N (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_RESET_B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_SCE (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SCD (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_Y (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_RESET_B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_D (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_D_N (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_SCE (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_RESET_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_Y (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net238_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_Y (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_S0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_Y (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_SCD (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_SCD (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_SCE (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_Q_N (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_D (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SCD (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_Q (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_X (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A3 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_Q (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_X (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_C (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_Y (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A0 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_C1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A_N (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_X (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_D (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_SCD (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_S0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_DE (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_SET_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_X (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold20_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_B1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_SCE (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_Q_N (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold19_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_Q (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A_N (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_DE (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Q (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_SCD (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_SCD (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_RESET_B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_D (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_SET_B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_Y (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_D_N (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_SCE (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SET_B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SCD (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_SET_B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SCD (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_DE (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_SCD (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold12_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_A3 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A_N (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_Q (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_C (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCE (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_Q (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_RESET_B (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_SCD (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_SCE (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCD (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_D (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_SCD (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_Y (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A_N (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_C (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_C (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_X (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_s763_GATE (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_X (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_Q (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_X (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_S0 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A3 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A_N (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_D1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_RESET_B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_Y (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A3 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_Q_N (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_RESET_B (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_B_N (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_Q (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_C_N (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_D (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_C_N (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_C (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_B1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_Y (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SCD (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_D (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_SCD (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCD (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SCD (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_Y (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_SCD (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_Q (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_Q_N (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCE (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_D1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_SCD (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCE (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_Q_N (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_SCD (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_Q (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_SCE (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_Q_N (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_B (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_Q (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A0 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_X (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_SCD (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_Q (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_C (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_X (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_RESET_B (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_SET_B (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_X (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_RESET_B (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_Q (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_B (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_SCD (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c642_Q (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_D (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_C1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_RESET_B (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A3 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_Q (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_C (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SCD (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_Q (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_B1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_SCE (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_Q (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_D1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_X (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold26_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_s750_Q_N (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_D1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone9_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold54_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_s777_Q (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SET_B (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SET_B (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_D1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_B_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_D1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_D_N (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_s804_Q (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_D1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A_N (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B_N (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_C1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A_N (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_D_N (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_Y (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_RESET_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_D1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_C1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_D1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_C (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_Y (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B_N (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_D_N (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_Y (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A_N (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_D1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_D1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A_N (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_B (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_C_N (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_C_N (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_B (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone9_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_C1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B_N (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A0 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A_N (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_D (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_S0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_B (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_D (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_S1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_C (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_A_N (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_C (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A_N (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_RESET_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A_N (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_C1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_RESET_B (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_C (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_RESET_B (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_C_N (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_C_N (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_D (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_S1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_C (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A_N (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_C_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_D_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_C_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_C1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_C (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_C1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_C (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_C_N (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A_N (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_C_N (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B_N (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_C1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_A_N (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A_N (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_D (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net794_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_SCE (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_s798_Q (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_s755_Q (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net801_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_Y (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_B (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_Q (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_s750_Q (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A3 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_D1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_C_N (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_Q (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net815_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_s802_Q (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_D_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_C (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_SCE (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_RESET_B (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B_N (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_Q (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_C_N (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_Y (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_C_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_Y (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap124_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_SCD (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_B_N (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire125_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SCD (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_SCE (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_SCE (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_C (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_D_N (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_C_N (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_SET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_C_N (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap133_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap137_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_C (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_C_N (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_D1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_SCE (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_B1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_D1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_SET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_D_N (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_B1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_C (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_C (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_D1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_D1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_SCD (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire144_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_D (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_C_N (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_RESET_B (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_C_N (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_D1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_B (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_D1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_S1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_C1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_C1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_D1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_D (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_SCE (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap149_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire148_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_D1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_C1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_C (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_C (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_C (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_D_N (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B_N (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_S0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_C (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_SCE (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C_N (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SET_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_SET_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SCE (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_RESET_B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_SCE (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_D_N (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_D1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_C (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_D1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_C1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_C_N (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_C1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_S0 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A0 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCD (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_SCD (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net476_X (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_RESET_B (.DIODE(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net476_X (.DIODE(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_S1 (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_C1 (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_SCE (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net671_X (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_C1 (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_D (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net794_X (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_RESET_B (.DIODE(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net238_X (.DIODE(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SET_B (.DIODE(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCE (.DIODE(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net238_X (.DIODE(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A1 (.DIODE(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net815_X (.DIODE(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_C (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_C (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_SET_B (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_RESET_B (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net843_X (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net379_X (.DIODE(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_SCD (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_C1 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_D (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net142_X (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_D_N (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_D1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_D_N (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_C (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_C (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_D_N (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net142_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net818_X (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_SCD (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S1 (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net818_X (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_RESET_B (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net801_X (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net801_X (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_C (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_B1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_D (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_Y (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_D_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_D1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_SCD (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_SET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone7_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone9_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net755));
 sky130_fd_sc_hd__mux4_1 clone2 (.A0(net739),
    .A1(net733),
    .A2(net743),
    .A3(net735),
    .S0(net63),
    .S1(net895),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net365),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net964),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net964),
    .X(net966));
 sky130_fd_sc_hd__and2_1 clone10 (.A(net16),
    .B(net732),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer12 (.A(net139),
    .X(net968));
 sky130_fd_sc_hd__and3_1 clone13 (.A(net970),
    .B(net742),
    .C(net734),
    .X(net969));
 sky130_fd_sc_hd__mux4_1 clone14 (.A0(net739),
    .A1(net733),
    .A2(net743),
    .A3(net735),
    .S0(net63),
    .S1(net895),
    .X(net970));
 sky130_fd_sc_hd__and2b_1 clone15 (.A_N(net87),
    .B(net78),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_1 rebuffer16 (.A(net13),
    .X(net972));
 sky130_fd_sc_hd__nand2_1 clone17 (.A(net4),
    .B(net3),
    .Y(net973));
 sky130_fd_sc_hd__clkbuf_1 clone18 (.A(in7),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(clknet_0_net142),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(clknet_0_net142),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_1 rebuffer21 (.A(clknet_1_0__leaf_net145),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(clknet_1_0__leaf_net145),
    .X(net978));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
