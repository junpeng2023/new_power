module netlist_1 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input in52,
	input in53,
	input in54,
	input in55,
	input in56,
	input in57,
	input in58,
	input in59,
	input in60,
	input in61,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51,
	output out52,
	output out53,
	output out54,
	output out55,
	output out56,
	output out57,
	output out58,
	output out59,
	output out60,
	output out61
);


wire net669;
wire net668;
wire net667;
wire net664;
wire net659;
wire net656;
wire out30;
wire net652;
wire net651;
wire net645;
wire net641;
wire net637;
wire net632;
wire net631;
wire net629;
wire net628;
wire net627;
wire net626;
wire net624;
wire net623;
wire net620;
wire net619;
wire net615;
wire net614;
wire net613;
wire net612;
wire net638;
wire net610;
wire net608;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire net596;
wire net592;
wire net588;
wire net587;
wire net583;
wire net582;
wire net584;
wire net581;
wire net579;
wire net577;
wire net576;
wire net569;
wire net567;
wire net566;
wire net565;
wire net562;
wire net559;
wire net556;
wire net647;
wire net555;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire net550;
wire net544;
wire net539;
wire net534;
wire net532;
wire net530;
wire net617;
wire net537;
wire net528;
wire net525;
wire net523;
wire net520;
wire net519;
wire net516;
wire net514;
wire net508;
wire net504;
wire net503;
wire net499;
wire clk;
wire net496;
wire net495;
wire net494;
wire net493;
wire net492;
wire net491;
wire net490;
wire net489;
wire net487;
wire net486;
wire out20;
wire net478;
wire net474;
wire net473;
wire net472;
wire net468;
wire net540;
wire net465;
wire net462;
wire net469;
wire net461;
wire net546;
wire net460;
wire net454;
wire net453;
wire net648;
wire net452;
wire net449;
wire net448;
wire net498;
wire net446;
wire net444;
wire out7;
wire net442;
wire out15;
wire net441;
wire net609;
wire net440;
wire net439;
wire net438;
wire net433;
wire net432;
wire net431;
wire net430;
wire net618;
wire net429;
wire net428;
wire net427;
wire net426;
wire net425;
wire net423;
wire net531;
wire net421;
wire net420;
wire net450;
wire net418;
wire net415;
wire net414;
wire net413;
wire net412;
wire net411;
wire net410;
wire net409;
wire net407;
wire out19;
wire net406;
wire net662;
wire net405;
wire net607;
wire net526;
wire net404;
wire net403;
wire net663;
wire net402;
wire net572;
wire net401;
wire net399;
wire net398;
wire net476;
wire net396;
wire net391;
wire net557;
wire net527;
wire net488;
wire net390;
wire net646;
wire net389;
wire net513;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net380;
wire net379;
wire net616;
wire net378;
wire net377;
wire net376;
wire out21;
wire net625;
wire net598;
wire net374;
wire out13;
wire net373;
wire net372;
wire net371;
wire net370;
wire net368;
wire net367;
wire net366;
wire net365;
wire net364;
wire net363;
wire net360;
wire net397;
wire net357;
wire net356;
wire net355;
wire out17;
wire net590;
wire net507;
wire net351;
wire net350;
wire net547;
wire net511;
wire net343;
wire net666;
wire net340;
wire net339;
wire net337;
wire net336;
wire net538;
wire net334;
wire net333;
wire net332;
wire net331;
wire net517;
wire net328;
wire net327;
wire out43;
wire net325;
wire net324;
wire net321;
wire net535;
wire net320;
wire net318;
wire net315;
wire net313;
wire net505;
wire net319;
wire net312;
wire out14;
wire net309;
wire net308;
wire net352;
wire net307;
wire net305;
wire net303;
wire net417;
wire out8;
wire net302;
wire net301;
wire net298;
wire net463;
wire net297;
wire net296;
wire net293;
wire in4;
wire out39;
wire net292;
wire net500;
wire net445;
wire out22;
wire net291;
wire net665;
wire net422;
wire net289;
wire net482;
wire in25;
wire net288;
wire net589;
wire net424;
wire net278;
wire net276;
wire net274;
wire net643;
wire net273;
wire out10;
wire in39;
wire net272;
wire net114;
wire net270;
wire in17;
wire net267;
wire net644;
wire net266;
wire out27;
wire net475;
wire net102;
wire net151;
wire net264;
wire net657;
wire net591;
wire net262;
wire net217;
wire net261;
wire net153;
wire out61;
wire net316;
wire out31;
wire net257;
wire net117;
wire net62;
wire net254;
wire net203;
wire net253;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire net661;
wire net241;
wire out42;
wire net238;
wire net142;
wire net183;
wire net234;
wire net232;
wire out12;
wire net226;
wire net524;
wire net382;
wire net259;
wire net335;
wire net222;
wire net219;
wire net578;
wire net210;
wire net213;
wire net208;
wire out16;
wire net188;
wire net207;
wire out56;
wire out38;
wire net649;
wire net205;
wire net202;
wire net199;
wire net384;
wire net224;
wire net122;
wire net197;
wire net193;
wire net192;
wire net190;
wire in20;
wire net189;
wire net246;
wire net186;
wire net126;
wire net284;
wire net655;
wire net563;
wire net549;
wire net182;
wire net342;
wire net17;
wire out44;
wire net310;
wire in49;
wire net147;
wire net180;
wire out23;
wire out40;
wire net258;
wire net464;
wire net3;
wire net176;
wire net133;
wire net175;
wire net573;
wire net240;
wire net416;
wire out33;
wire net173;
wire net595;
wire out52;
wire net195;
wire net479;
wire net8;
wire net172;
wire net622;
wire net518;
wire net170;
wire net381;
wire net218;
wire net169;
wire net344;
wire net168;
wire net286;
wire net167;
wire net58;
wire net221;
wire net166;
wire net269;
wire net165;
wire net660;
wire net359;
wire out28;
wire out60;
wire out45;
wire net497;
wire net161;
wire net285;
wire net160;
wire net636;
wire net311;
wire in37;
wire net159;
wire net158;
wire out58;
wire out6;
wire net152;
wire net150;
wire net149;
wire net148;
wire net178;
wire net239;
wire net144;
wire net322;
wire net299;
wire net143;
wire out37;
wire out57;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net561;
wire out29;
wire net139;
wire net137;
wire net136;
wire net456;
wire net135;
wire net157;
wire net177;
wire out51;
wire net134;
wire net250;
wire net225;
wire net132;
wire net201;
wire net130;
wire net358;
wire net294;
wire net127;
wire net124;
wire net640;
wire net369;
wire net50;
wire out18;
wire net255;
wire net548;
wire net481;
wire net383;
wire net120;
wire net204;
wire out0;
wire net164;
wire net110;
wire net109;
wire net642;
wire net268;
wire in7;
wire net82;
wire net123;
wire net282;
wire net71;
wire net229;
wire net326;
wire net108;
wire net107;
wire net104;
wire in12;
wire net271;
wire net103;
wire net408;
wire out26;
wire net99;
wire net6;
wire out50;
wire net348;
wire net341;
wire in52;
wire net96;
wire net466;
wire net118;
wire net94;
wire net90;
wire net74;
wire net277;
wire net639;
wire net88;
wire net81;
wire net230;
wire net156;
wire net361;
wire net115;
wire net670;
wire net209;
wire in18;
wire net34;
wire net79;
wire net231;
wire net349;
wire net329;
wire net212;
wire net653;
wire net485;
wire net78;
wire in5;
wire net77;
wire net76;
wire net236;
wire net571;
wire net31;
wire net73;
wire net116;
wire net69;
wire net128;
wire net67;
wire net447;
wire net98;
wire net522;
wire net459;
wire net436;
wire out9;
wire net260;
wire net541;
wire net501;
wire net323;
wire net15;
wire net64;
wire net63;
wire net354;
wire in38;
wire net198;
wire net467;
wire net101;
wire net9;
wire net306;
wire net75;
wire in56;
wire out48;
wire net61;
wire net512;
wire out34;
wire net179;
wire net60;
wire net237;
wire net59;
wire net248;
wire net275;
wire net119;
wire net477;
wire net400;
wire in10;
wire net228;
wire net39;
wire net630;
wire net56;
wire out53;
wire net55;
wire net244;
wire net568;
wire net223;
wire net330;
wire out32;
wire net214;
wire net53;
wire net97;
wire in48;
wire net196;
wire net52;
wire net597;
wire out55;
wire net155;
wire net338;
wire net46;
wire in31;
wire net65;
wire net392;
wire net113;
wire net575;
wire net434;
wire net200;
wire net162;
wire net395;
wire out3;
wire net564;
wire net443;
wire net154;
wire net345;
wire net84;
wire in46;
wire net85;
wire net72;
wire net131;
wire net502;
wire net235;
wire net49;
wire net594;
wire net215;
wire net484;
wire net184;
wire in8;
wire net346;
wire net43;
wire net599;
wire net112;
wire net650;
wire net185;
wire net585;
wire net560;
wire net45;
wire net252;
wire net38;
wire net187;
wire in13;
wire net621;
wire net586;
wire net533;
wire net32;
wire net419;
wire net125;
wire net458;
wire net19;
wire net347;
wire in15;
wire net20;
wire in19;
wire net27;
wire net70;
wire net48;
wire net28;
wire net92;
wire net25;
wire net30;
wire net29;
wire net570;
wire out2;
wire in0;
wire net24;
wire out47;
wire net290;
wire net227;
wire out5;
wire net14;
wire out59;
wire net470;
wire net44;
wire net471;
wire in33;
wire net33;
wire net233;
wire net40;
wire in60;
wire net435;
wire net18;
wire net26;
wire net483;
wire net16;
wire net558;
wire in1;
wire net265;
wire net13;
wire net22;
wire net263;
wire net521;
wire net353;
wire out25;
wire out41;
wire net5;
wire net206;
wire in59;
wire in58;
wire net295;
wire in24;
wire in61;
wire net171;
wire in23;
wire in55;
wire out4;
wire net457;
wire net42;
wire net91;
wire net580;
wire net375;
wire in57;
wire net281;
wire net54;
wire net1;
wire in54;
wire in53;
wire out11;
wire net41;
wire net138;
wire net211;
wire in6;
wire net0;
wire in35;
wire net106;
wire in34;
wire net593;
wire in45;
wire net163;
wire net393;
wire net4;
wire in42;
wire net256;
wire net87;
wire net509;
wire net506;
wire net181;
wire net451;
wire net7;
wire out54;
wire out1;
wire net145;
wire net574;
wire net23;
wire net216;
wire net455;
wire net129;
wire net100;
wire net2;
wire in28;
wire in44;
wire net601;
wire out35;
wire in32;
wire in50;
wire net47;
wire net12;
wire in27;
wire in9;
wire net654;
wire net611;
wire net515;
wire net362;
wire in16;
wire net191;
wire out46;
wire net89;
wire in41;
wire in26;
wire net35;
wire net21;
wire net543;
wire net220;
wire in43;
wire net174;
wire in22;
wire net600;
wire net510;
wire net68;
wire in14;
wire net529;
wire in21;
wire net57;
wire net480;
wire net86;
wire net317;
wire in51;
wire net93;
wire net280;
wire in47;
wire in2;
wire net658;
wire net105;
wire in11;
wire net51;
wire net437;
wire in36;
wire net111;
wire net242;
wire net536;
wire net37;
wire net36;
wire net95;
wire net304;
wire net121;
wire net300;
wire in30;
wire net146;
wire net279;
wire net251;
wire net11;
wire net394;
wire net314;
wire in3;
wire net633;
wire net194;
wire net542;
wire net80;
wire in29;
sky130_fd_sc_hd__mux4_2 c62(
.A0(in49),
.A1(in23),
.A2(in60),
.A3(in61),
.S0(in39),
.S1(net3),
.X(net0)
);

sky130_fd_sc_hd__mux4_2 c63(
.A0(in53),
.A1(in57),
.A2(in39),
.A3(in56),
.S0(in3),
.S1(in61),
.X(net1)
);

sky130_fd_sc_hd__mux4_1 c64(
.A0(in38),
.A1(in44),
.A2(in59),
.A3(in46),
.S0(in45),
.S1(in58),
.X(net2)
);

sky130_fd_sc_hd__a211oi_4 c65(
.A1(in3),
.A2(in28),
.B1(in39),
.C1(in14),
.Y(net3)
);

sky130_fd_sc_hd__or2_4 c66(
.A(in45),
.B(in47),
.X(net4)
);

sky130_fd_sc_hd__nor2b_1 c67(
.A(in32),
.B_N(in50),
.Y(net5)
);

sky130_fd_sc_hd__and2_4 c68(
.A(in61),
.B(in53),
.X(net6)
);

sky130_fd_sc_hd__or2b_4 c69(
.A(net5),
.B_N(in23),
.X(net7)
);

sky130_fd_sc_hd__nor2_4 c70(
.A(net7),
.B(in45),
.Y(net8)
);

sky130_fd_sc_hd__and2_4 c71(
.A(in49),
.B(net8),
.X(net9)
);

sky130_fd_sc_hd__nor2b_4 c72(
.A(in60),
.B_N(in11),
.Y(net10)
);

sky130_fd_sc_hd__and2_0 c73(
.A(in34),
.B(net10),
.X(net11)
);

sky130_fd_sc_hd__and2_2 c74(
.A(net1),
.B(in23),
.X(net12)
);

sky130_fd_sc_hd__and2_2 c75(
.A(in23),
.B(net11),
.X(net13)
);

sky130_fd_sc_hd__and2_2 c76(
.A(net10),
.B(net12),
.X(net14)
);

sky130_fd_sc_hd__nor3_1 c77(
.A(net11),
.B(net1),
.C(net12),
.Y(net15)
);

sky130_fd_sc_hd__and2b_4 c78(
.A_N(net13),
.B(net15),
.X(net16)
);

sky130_fd_sc_hd__and3b_4 c79(
.A_N(net15),
.B(net13),
.C(in45),
.X(net17)
);

sky130_fd_sc_hd__and2b_4 c80(
.A_N(net12),
.B(net17),
.X(net18)
);

sky130_fd_sc_hd__and2b_4 c81(
.A_N(net18),
.B(net12),
.X(net19)
);

sky130_fd_sc_hd__mux4_1 c82(
.A0(in56),
.A1(net18),
.A2(net19),
.A3(net13),
.S0(net11),
.S1(net9),
.X(net20)
);

sky130_fd_sc_hd__or3_4 c83(
.A(in40),
.B(net13),
.C(net19),
.X(net21)
);

sky130_fd_sc_hd__nand3_1 c84(
.A(net21),
.B(net6),
.C(net18),
.Y(net22)
);

sky130_fd_sc_hd__mux4_1 c85(
.A0(in33),
.A1(net22),
.A2(net12),
.A3(net18),
.S0(net13),
.S1(net5),
.X(out25)
);

sky130_fd_sc_hd__nor3_2 c86(
.A(net20),
.B(net9),
.C(net22),
.Y(net23)
);

sky130_fd_sc_hd__nor3b_1 c87(
.A(net14),
.B(net11),
.C_N(net23),
.Y(net24)
);

sky130_fd_sc_hd__or2_2 c88(
.A(in53),
.B(net19),
.X(net25)
);

sky130_fd_sc_hd__nand2b_4 c89(
.A_N(net20),
.B(in7),
.Y(net26)
);

sky130_fd_sc_hd__and2_1 c90(
.A(net17),
.B(in53),
.X(net27)
);

sky130_fd_sc_hd__and2b_2 c91(
.A_N(net26),
.B(net27),
.X(net28)
);

sky130_fd_sc_hd__or2b_1 c92(
.A(net26),
.B_N(in21),
.X(net29)
);

sky130_fd_sc_hd__or2b_4 c93(
.A(net29),
.B_N(net24),
.X(net30)
);

sky130_fd_sc_hd__nand2_1 c94(
.A(net19),
.B(in7),
.Y(net31)
);

sky130_fd_sc_hd__a211o_1 c95(
.A1(net8),
.A2(net27),
.B1(net26),
.C1(in55),
.X(net32)
);

sky130_fd_sc_hd__nor2_4 c96(
.A(net13),
.B(net29),
.Y(net33)
);

sky130_fd_sc_hd__or2_2 c97(
.A(net32),
.B(net30),
.X(net34)
);

sky130_fd_sc_hd__nor2_4 c98(
.A(net34),
.B(net16),
.Y(net35)
);

sky130_fd_sc_hd__nor2b_1 c99(
.A(net6),
.B_N(net28),
.Y(net36)
);

sky130_fd_sc_hd__nand2_1 c100(
.A(net22),
.B(net29),
.Y(out22)
);

sky130_fd_sc_hd__or2b_4 c101(
.A(in39),
.B_N(net29),
.X(net37)
);

sky130_fd_sc_hd__nor2_4 c102(
.A(out22),
.B(net14),
.Y(net38)
);

sky130_fd_sc_hd__nand2b_2 c103(
.A_N(net37),
.B(net25),
.Y(net39)
);

sky130_fd_sc_hd__or2b_4 c104(
.A(net35),
.B_N(net8),
.X(out16)
);

sky130_fd_sc_hd__or2b_4 c105(
.A(net25),
.B_N(net39),
.X(net40)
);

sky130_fd_sc_hd__and2_2 c106(
.A(net36),
.B(net40),
.X(net41)
);

sky130_fd_sc_hd__a211o_2 c107(
.A1(net35),
.A2(net31),
.B1(out22),
.C1(net29),
.X(net42)
);

sky130_fd_sc_hd__a211oi_4 c108(
.A1(net40),
.A2(net41),
.B1(net37),
.C1(net42),
.Y(net43)
);

sky130_fd_sc_hd__mux4_4 c109(
.A0(net42),
.A1(net25),
.A2(net40),
.A3(net41),
.S0(net43),
.S1(net29),
.X(net44)
);

sky130_fd_sc_hd__dfbbn_1 c110(
.D(net43),
.RESET_B(net39),
.SET_B(net28),
.CLK_N(clk),
.Q(out57),
.Q_N(net45)
);

sky130_fd_sc_hd__or2_1 c111(
.A(net29),
.B(in26),
.X(out3)
);

sky130_fd_sc_hd__and2_1 c112(
.A(in50),
.B(net29),
.X(out53)
);

sky130_fd_sc_hd__nand3_2 c113(
.A(net36),
.B(out57),
.C(net12),
.Y(net46)
);

sky130_fd_sc_hd__nor2_1 c114(
.A(net12),
.B(net36),
.Y(net47)
);

sky130_fd_sc_hd__and2b_4 c115(
.A_N(in61),
.B(net652),
.X(net48)
);

sky130_fd_sc_hd__nand2b_2 c116(
.A_N(net39),
.B(in61),
.Y(net49)
);

sky130_fd_sc_hd__and3b_2 c117(
.A_N(net15),
.B(in61),
.C(net47),
.X(net50)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c118(
.A(net636),
.X(net51)
);

sky130_fd_sc_hd__nor2b_1 c119(
.A(net24),
.B_N(net49),
.Y(net52)
);

sky130_fd_sc_hd__nor3b_2 c120(
.A(net51),
.B(out16),
.C_N(out22),
.Y(net53)
);

sky130_fd_sc_hd__or2_2 c121(
.A(net47),
.B(net28),
.X(out32)
);

sky130_fd_sc_hd__buf_1 c122(
.A(net636),
.X(net54)
);

sky130_fd_sc_hd__a211o_2 c123(
.A1(out32),
.A2(net45),
.B1(out3),
.C1(in26),
.X(net55)
);

sky130_fd_sc_hd__dfbbn_2 c124(
.D(net53),
.RESET_B(net49),
.SET_B(net36),
.CLK_N(clk),
.Q(net57),
.Q_N(net56)
);

sky130_fd_sc_hd__dfbbp_1 c125(
.D(net49),
.RESET_B(net56),
.SET_B(net53),
.CLK(clk),
.Q(net59),
.Q_N(net58)
);

sky130_fd_sc_hd__mux4_4 c126(
.A0(net28),
.A1(net49),
.A2(net58),
.A3(net43),
.S0(out16),
.S1(in61),
.X(net60)
);

sky130_fd_sc_hd__sdfxbp_1 c127(
.D(net57),
.SCD(net58),
.SCE(net53),
.CLK(clk),
.Q(out48),
.Q_N(net61)
);

sky130_fd_sc_hd__a211o_1 c128(
.A1(net59),
.A2(net21),
.B1(net54),
.C1(net653),
.X(out51)
);

sky130_fd_sc_hd__sdfrbp_1 c129(
.D(out51),
.RESET_B(out16),
.SCD(net43),
.SCE(net654),
.CLK(clk),
.Q(net62)
);

sky130_fd_sc_hd__and3b_1 c130(
.A_N(net62),
.B(net49),
.C(out51),
.X(out47)
);

sky130_fd_sc_hd__and3_1 c131(
.A(net51),
.B(net59),
.C(out51),
.X(net63)
);

sky130_fd_sc_hd__and2b_1 c132(
.A_N(in9),
.B(in10),
.X(net64)
);

sky130_fd_sc_hd__nor2_4 c133(
.A(net64),
.B(in15),
.Y(net65)
);

sky130_fd_sc_hd__nor2b_2 c134(
.A(in18),
.B_N(in2),
.Y(net66)
);

sky130_fd_sc_hd__nand2_2 c135(
.A(in2),
.B(in18),
.Y(net67)
);

sky130_fd_sc_hd__or2_1 c136(
.A(net65),
.B(in17),
.X(net68)
);

sky130_fd_sc_hd__nand2_2 c137(
.A(net65),
.B(net66),
.Y(net69)
);

sky130_fd_sc_hd__nor2b_2 c138(
.A(in13),
.B_N(in21),
.Y(net70)
);

sky130_fd_sc_hd__nor2b_1 c139(
.A(net69),
.B_N(in20),
.Y(net71)
);

sky130_fd_sc_hd__and2_4 c140(
.A(net68),
.B(net71),
.X(net72)
);

sky130_fd_sc_hd__or2b_4 c141(
.A(net70),
.B_N(in19),
.X(net73)
);

sky130_fd_sc_hd__and2b_4 c142(
.A_N(net65),
.B(net69),
.X(net74)
);

sky130_fd_sc_hd__nor2_2 c143(
.A(in15),
.B(net73),
.Y(net75)
);

sky130_fd_sc_hd__a211o_1 c144(
.A1(in19),
.A2(in5),
.B1(in20),
.C1(in13),
.X(net76)
);

sky130_fd_sc_hd__nand3b_4 c145(
.A_N(net76),
.B(net75),
.C(net71),
.Y(net77)
);

sky130_fd_sc_hd__or2_1 c146(
.A(net67),
.B(net75),
.X(net78)
);

sky130_fd_sc_hd__or3_4 c147(
.A(net78),
.B(net77),
.C(net76),
.X(net79)
);

sky130_fd_sc_hd__nor2b_4 c148(
.A(net75),
.B_N(net74),
.Y(net80)
);

sky130_fd_sc_hd__and2b_2 c149(
.A_N(net66),
.B(net76),
.X(net81)
);

sky130_fd_sc_hd__nand2b_1 c150(
.A_N(net80),
.B(net81),
.Y(net82)
);

sky130_fd_sc_hd__mux4_4 c151(
.A0(net75),
.A1(net79),
.A2(in18),
.A3(net78),
.S0(in9),
.S1(in15),
.X(net83)
);

sky130_fd_sc_hd__and3b_1 c152(
.A_N(net72),
.B(net74),
.C(net81),
.X(net84)
);

sky130_fd_sc_hd__a311oi_2 c153(
.A1(net84),
.A2(net71),
.A3(net83),
.B1(net79),
.C1(net72),
.Y(net85)
);

sky130_fd_sc_hd__or2_4 c154(
.A(net82),
.B(in16),
.X(net86)
);

sky130_fd_sc_hd__and2b_2 c155(
.A_N(in12),
.B(in14),
.X(net87)
);

sky130_fd_sc_hd__and2b_1 c156(
.A_N(net87),
.B(in22),
.X(net88)
);

sky130_fd_sc_hd__or3b_1 c157(
.A(net88),
.B(in28),
.C_N(in29),
.X(net89)
);

sky130_fd_sc_hd__nand2b_1 c158(
.A_N(in29),
.B(in24),
.Y(net90)
);

sky130_fd_sc_hd__nor3_2 c159(
.A(net90),
.B(in27),
.C(net86),
.Y(net91)
);

sky130_fd_sc_hd__nand2_2 c160(
.A(in16),
.B(net78),
.Y(net92)
);

sky130_fd_sc_hd__nand2_2 c161(
.A(in36),
.B(net87),
.Y(net93)
);

sky130_fd_sc_hd__nand2b_1 c162(
.A_N(in24),
.B(in29),
.Y(net94)
);

sky130_fd_sc_hd__nand2_1 c163(
.A(net77),
.B(net88),
.Y(net95)
);

sky130_fd_sc_hd__or3b_4 c164(
.A(net85),
.B(in10),
.C_N(net93),
.X(net96)
);

sky130_fd_sc_hd__nor2b_2 c165(
.A(net73),
.B_N(net90),
.Y(net97)
);

sky130_fd_sc_hd__nand2_2 c166(
.A(net97),
.B(in24),
.Y(net98)
);

sky130_fd_sc_hd__or2_2 c167(
.A(in41),
.B(net94),
.X(net99)
);

sky130_fd_sc_hd__a211o_2 c168(
.A1(in31),
.A2(net85),
.B1(net81),
.C1(net97),
.X(net100)
);

sky130_fd_sc_hd__and2_4 c169(
.A(net79),
.B(net99),
.X(net101)
);

sky130_fd_sc_hd__and2_0 c170(
.A(net101),
.B(net82),
.X(net102)
);

sky130_fd_sc_hd__mux4_2 c171(
.A0(in42),
.A1(net91),
.A2(net100),
.A3(net96),
.S0(in7),
.S1(in28),
.X(net103)
);

sky130_fd_sc_hd__a311oi_1 c172(
.A1(net92),
.A2(net87),
.A3(net102),
.B1(net101),
.C1(net97),
.Y(net104)
);

sky130_fd_sc_hd__and3_1 c173(
.A(net70),
.B(net104),
.C(net97),
.X(net105)
);

sky130_fd_sc_hd__nand3b_1 c174(
.A_N(net100),
.B(net104),
.C(net78),
.Y(net106)
);

sky130_fd_sc_hd__nand3_2 c175(
.A(net106),
.B(net105),
.C(net104),
.Y(net107)
);

sky130_fd_sc_hd__and2_2 c176(
.A(net81),
.B(net96),
.X(net108)
);

sky130_fd_sc_hd__nor2b_4 c177(
.A(net104),
.B_N(net3),
.Y(net109)
);

sky130_fd_sc_hd__nand3b_1 c178(
.A_N(net86),
.B(net89),
.C(in48),
.Y(net110)
);

sky130_fd_sc_hd__nor2b_4 c179(
.A(in30),
.B_N(net93),
.Y(net111)
);

sky130_fd_sc_hd__and2b_1 c180(
.A_N(net96),
.B(in44),
.X(net112)
);

sky130_fd_sc_hd__nand2_2 c181(
.A(in59),
.B(net84),
.Y(net113)
);

sky130_fd_sc_hd__nand2b_2 c182(
.A_N(in43),
.B(net109),
.Y(net114)
);

sky130_fd_sc_hd__nand2_4 c183(
.A(in46),
.B(net103),
.Y(net115)
);

sky130_fd_sc_hd__or2_4 c184(
.A(net3),
.B(net109),
.X(net116)
);

sky130_fd_sc_hd__and2b_2 c185(
.A_N(in22),
.B(net3),
.X(net117)
);

sky130_fd_sc_hd__nand2_2 c186(
.A(net114),
.B(in51),
.Y(net118)
);

sky130_fd_sc_hd__nand2b_2 c187(
.A_N(net0),
.B(net118),
.Y(net119)
);

sky130_fd_sc_hd__nand2b_1 c188(
.A_N(net111),
.B(net3),
.Y(net120)
);

sky130_fd_sc_hd__nand2b_4 c189(
.A_N(net110),
.B(in25),
.Y(net121)
);

sky130_fd_sc_hd__and2b_4 c190(
.A_N(net109),
.B(in57),
.X(out12)
);

sky130_fd_sc_hd__or3b_1 c191(
.A(net117),
.B(net121),
.C_N(out12),
.X(net122)
);

sky130_fd_sc_hd__and2b_4 c192(
.A_N(net118),
.B(out12),
.X(net123)
);

sky130_fd_sc_hd__or3b_2 c193(
.A(net116),
.B(net112),
.C_N(in28),
.X(net124)
);

sky130_fd_sc_hd__a211o_4 c194(
.A1(net115),
.A2(net112),
.B1(net118),
.C1(out12),
.X(net125)
);

sky130_fd_sc_hd__or2_1 c195(
.A(net122),
.B(out12),
.X(net126)
);

sky130_fd_sc_hd__or3b_4 c196(
.A(net126),
.B(net115),
.C_N(net117),
.X(net127)
);

sky130_fd_sc_hd__nor2_2 c197(
.A(net123),
.B(net126),
.Y(net128)
);

sky130_fd_sc_hd__nand2_4 c198(
.A(in51),
.B(net128),
.Y(net129)
);

sky130_fd_sc_hd__sdfxbp_2 c199(
.D(in58),
.SCD(in27),
.SCE(net129),
.CLK(clk),
.Q(net130)
);

sky130_fd_sc_hd__or2_2 c200(
.A(net128),
.B(in48),
.X(net131)
);

sky130_fd_sc_hd__or2_4 c201(
.A(net99),
.B(net125),
.X(net132)
);

sky130_fd_sc_hd__buf_16 c202(
.A(net617),
.X(net133)
);

sky130_fd_sc_hd__or2b_4 c203(
.A(net4),
.B_N(net113),
.X(net134)
);

sky130_fd_sc_hd__and2b_1 c204(
.A_N(net89),
.B(in51),
.X(net135)
);

sky130_fd_sc_hd__clkinv_4 c205(
.A(net616),
.Y(net136)
);

sky130_fd_sc_hd__nor2_2 c206(
.A(net117),
.B(net67),
.Y(net137)
);

sky130_fd_sc_hd__and2_4 c207(
.A(net130),
.B(net119),
.X(net138)
);

sky130_fd_sc_hd__nor2_1 c208(
.A(net136),
.B(net134),
.Y(net139)
);

sky130_fd_sc_hd__clkinv_16 c209(
.A(net651),
.Y(net140)
);

sky130_fd_sc_hd__and2_1 c210(
.A(net138),
.B(in27),
.X(net141)
);

sky130_fd_sc_hd__clkinv_1 c211(
.A(net651),
.Y(net142)
);

sky130_fd_sc_hd__dfrbp_1 c212(
.D(net125),
.RESET_B(net131),
.CLK(clk),
.Q(net144),
.Q_N(net143)
);

sky130_fd_sc_hd__inv_12 c213(
.A(net650),
.Y(net145)
);

sky130_fd_sc_hd__nand3_1 c214(
.A(in52),
.B(net99),
.C(net145),
.Y(net146)
);

sky130_fd_sc_hd__nor2_4 c215(
.A(net120),
.B(out12),
.Y(net147)
);

sky130_fd_sc_hd__or2_4 c216(
.A(net147),
.B(net142),
.X(net148)
);

sky130_fd_sc_hd__or3_1 c217(
.A(net132),
.B(net135),
.C(net4),
.X(net149)
);

sky130_fd_sc_hd__nand3_1 c218(
.A(net146),
.B(net148),
.C(net147),
.Y(net150)
);

sky130_fd_sc_hd__nor3b_4 c219(
.A(net23),
.B(net150),
.C_N(net146),
.Y(net151)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c220(
.A(net612),
.X(net152)
);

sky130_fd_sc_hd__and2b_1 c221(
.A_N(net34),
.B(net145),
.X(out6)
);

sky130_fd_sc_hd__nand2_1 c222(
.A(out6),
.B(net103),
.Y(net153)
);

sky130_fd_sc_hd__inv_12 c223(
.A(net611),
.Y(net154)
);

sky130_fd_sc_hd__and3_1 c224(
.A(in54),
.B(net98),
.C(net34),
.X(net155)
);

sky130_fd_sc_hd__nand2_2 c225(
.A(net5),
.B(out6),
.Y(out58)
);

sky130_fd_sc_hd__nor3b_1 c226(
.A(net67),
.B(net2),
.C_N(net5),
.Y(net156)
);

sky130_fd_sc_hd__nor3_2 c227(
.A(net27),
.B(in27),
.C(net148),
.Y(net157)
);

sky130_fd_sc_hd__or2_2 c228(
.A(net137),
.B(out6),
.X(net158)
);

sky130_fd_sc_hd__or2b_1 c229(
.A(net155),
.B_N(net16),
.X(net159)
);

sky130_fd_sc_hd__or2_1 c230(
.A(net156),
.B(out58),
.X(out1)
);

sky130_fd_sc_hd__dfrbp_2 c231(
.D(net151),
.RESET_B(net38),
.CLK(clk),
.Q(net161),
.Q_N(net160)
);

sky130_fd_sc_hd__nor3b_1 c232(
.A(net156),
.B(out12),
.C_N(net16),
.Y(net162)
);

sky130_fd_sc_hd__or3b_2 c233(
.A(net161),
.B(net157),
.C_N(net67),
.X(out28)
);

sky130_fd_sc_hd__nor2_1 c234(
.A(net41),
.B(net145),
.Y(net163)
);

sky130_fd_sc_hd__mux4_1 c235(
.A0(net152),
.A1(net155),
.A2(net160),
.A3(in54),
.S0(net134),
.S1(net154),
.X(net164)
);

sky130_fd_sc_hd__nor2b_2 c236(
.A(net162),
.B_N(net163),
.Y(net165)
);

sky130_fd_sc_hd__dfrtn_1 c237(
.D(net98),
.RESET_B(out28),
.CLK_N(clk),
.Q(out11)
);

sky130_fd_sc_hd__sdfxtp_1 c238(
.D(net38),
.SCD(net161),
.SCE(out1),
.CLK(clk),
.Q(net166)
);

sky130_fd_sc_hd__a211o_2 c239(
.A1(net157),
.A2(out58),
.B1(net152),
.C1(net134),
.X(out46)
);

sky130_fd_sc_hd__sdfxtp_2 c240(
.D(net165),
.SCD(net98),
.SCE(out46),
.CLK(clk),
.Q(net167)
);

sky130_fd_sc_hd__mux4_2 c241(
.A0(net167),
.A1(net162),
.A2(out11),
.A3(net5),
.S0(net165),
.S1(net16),
.X(net168)
);

sky130_fd_sc_hd__nor2_2 c242(
.A(net31),
.B(out3),
.Y(net169)
);

sky130_fd_sc_hd__and2_4 c243(
.A(net48),
.B(net169),
.X(net170)
);

sky130_fd_sc_hd__or2_1 c244(
.A(net170),
.B(out25),
.X(net171)
);

sky130_fd_sc_hd__nand2_2 c245(
.A(net163),
.B(out25),
.Y(net172)
);

sky130_fd_sc_hd__or2_4 c246(
.A(net78),
.B(net652),
.X(out34)
);

sky130_fd_sc_hd__nand2b_2 c247(
.A_N(net54),
.B(net169),
.Y(net173)
);

sky130_fd_sc_hd__sdfbbn_1 c248(
.D(net154),
.RESET_B(out34),
.SCD(out22),
.SCE(net171),
.SET_B(net172),
.CLK_N(clk),
.Q(out33),
.Q_N(net174)
);

sky130_fd_sc_hd__inv_6 c249(
.A(net630),
.Y(net175)
);

sky130_fd_sc_hd__a211o_1 c250(
.A1(net55),
.A2(net61),
.B1(net78),
.C1(net45),
.X(net176)
);

sky130_fd_sc_hd__nand2_4 c251(
.A(net63),
.B(net48),
.Y(net177)
);

sky130_fd_sc_hd__nor2_4 c252(
.A(net177),
.B(net174),
.Y(net178)
);

sky130_fd_sc_hd__nor2_2 c253(
.A(net175),
.B(out34),
.Y(net179)
);

sky130_fd_sc_hd__nand2b_1 c254(
.A_N(net178),
.B(net179),
.Y(out59)
);

sky130_fd_sc_hd__sdfxtp_4 c255(
.D(net179),
.SCD(net172),
.SCE(out59),
.CLK(clk),
.Q(out54)
);

sky130_fd_sc_hd__nand2b_1 c256(
.A_N(net46),
.B(net178),
.Y(net180)
);

sky130_fd_sc_hd__a211o_4 c257(
.A1(net176),
.A2(net173),
.B1(out59),
.C1(net175),
.X(out42)
);

sky130_fd_sc_hd__or3b_1 c258(
.A(net169),
.B(net179),
.C_N(net180),
.X(out44)
);

sky130_fd_sc_hd__dlygate4sd1_1 c259(
.A(net629),
.X(out2)
);

sky130_fd_sc_hd__sdfbbn_2 c260(
.D(net178),
.RESET_B(out42),
.SCD(out22),
.SCE(out54),
.SET_B(net655),
.CLK_N(clk),
.Q(net181)
);

sky130_fd_sc_hd__dfbbn_1 c261(
.D(net158),
.RESET_B(out54),
.SET_B(out28),
.CLK_N(clk),
.Q(net183),
.Q_N(net182)
);

sky130_fd_sc_hd__or3_4 c262(
.A(net171),
.B(net183),
.C(in17),
.X(net184)
);

sky130_fd_sc_hd__a211oi_2 c263(
.A1(net184),
.A2(out2),
.B1(net171),
.C1(net182),
.Y(out40)
);

sky130_fd_sc_hd__and2b_4 c264(
.A_N(in8),
.B(net72),
.X(net185)
);

sky130_fd_sc_hd__and2_1 c265(
.A(in9),
.B(net84),
.X(net186)
);

sky130_fd_sc_hd__and2_0 c266(
.A(net68),
.B(net66),
.X(net187)
);

sky130_fd_sc_hd__nor2b_4 c267(
.A(net186),
.B_N(in12),
.Y(net188)
);

sky130_fd_sc_hd__nand3b_2 c268(
.A_N(net80),
.B(net187),
.C(net188),
.Y(net189)
);

sky130_fd_sc_hd__and2_2 c269(
.A(net185),
.B(net189),
.X(net190)
);

sky130_fd_sc_hd__nor2b_4 c270(
.A(net188),
.B_N(net189),
.Y(net191)
);

sky130_fd_sc_hd__nand2b_4 c271(
.A_N(in20),
.B(net83),
.Y(net192)
);

sky130_fd_sc_hd__nand2_2 c272(
.A(net192),
.B(net191),
.Y(net193)
);

sky130_fd_sc_hd__nand2_1 c273(
.A(net192),
.B(net193),
.Y(net194)
);

sky130_fd_sc_hd__or2_1 c274(
.A(net189),
.B(in14),
.X(net195)
);

sky130_fd_sc_hd__a311o_2 c275(
.A1(net195),
.A2(net74),
.A3(net185),
.B1(net193),
.C1(net187),
.X(net196)
);

sky130_fd_sc_hd__or2_2 c276(
.A(net72),
.B(net65),
.X(net197)
);

sky130_fd_sc_hd__or2b_4 c277(
.A(net186),
.B_N(net195),
.X(net198)
);

sky130_fd_sc_hd__nand2b_2 c278(
.A_N(net191),
.B(net66),
.Y(net199)
);

sky130_fd_sc_hd__and2b_2 c279(
.A_N(net199),
.B(net190),
.X(net200)
);

sky130_fd_sc_hd__nand2_4 c280(
.A(net194),
.B(net193),
.Y(net201)
);

sky130_fd_sc_hd__nand3b_2 c281(
.A_N(net201),
.B(net199),
.C(net187),
.Y(net202)
);

sky130_fd_sc_hd__nor2b_4 c282(
.A(net191),
.B_N(net200),
.Y(net203)
);

sky130_fd_sc_hd__nor3b_1 c283(
.A(net198),
.B(net187),
.C_N(net190),
.Y(net204)
);

sky130_fd_sc_hd__a211o_2 c284(
.A1(net202),
.A2(net201),
.B1(net186),
.C1(net188),
.X(net205)
);

sky130_fd_sc_hd__dlygate4sd1_1 c285(
.A(net649),
.X(out38)
);

sky130_fd_sc_hd__or2_1 c286(
.A(in35),
.B(in25),
.X(net206)
);

sky130_fd_sc_hd__or2_1 c287(
.A(in11),
.B(net197),
.X(net207)
);

sky130_fd_sc_hd__or2b_2 c288(
.A(in5),
.B_N(net206),
.X(out9)
);

sky130_fd_sc_hd__mux4_4 c289(
.A0(in37),
.A1(net84),
.A2(net92),
.A3(net65),
.S0(net97),
.S1(out9),
.X(net208)
);

sky130_fd_sc_hd__nor3_4 c290(
.A(net106),
.B(net107),
.C(in5),
.Y(net209)
);

sky130_fd_sc_hd__a21bo_1 c291(
.A1(net83),
.A2(net106),
.B1_N(net65),
.X(net210)
);

sky130_fd_sc_hd__a21oi_4 c292(
.A1(net206),
.A2(net93),
.B1(net208),
.Y(net211)
);

sky130_fd_sc_hd__nand2_4 c293(
.A(net210),
.B(net211),
.Y(net212)
);

sky130_fd_sc_hd__a21boi_4 c294(
.A1(net197),
.A2(net95),
.B1_N(net209),
.Y(net213)
);

sky130_fd_sc_hd__nor2b_2 c295(
.A(net213),
.B_N(in26),
.Y(net214)
);

sky130_fd_sc_hd__a21bo_1 c296(
.A1(net214),
.A2(net203),
.B1_N(out9),
.X(net215)
);

sky130_fd_sc_hd__nor2b_4 c297(
.A(net209),
.B_N(net105),
.Y(net216)
);

sky130_fd_sc_hd__a21o_1 c298(
.A1(net95),
.A2(out9),
.B1(net197),
.X(net217)
);

sky130_fd_sc_hd__o21ai_1 c299(
.A1(net212),
.A2(net217),
.B1(net209),
.Y(net218)
);

sky130_fd_sc_hd__and2b_1 c300(
.A_N(net107),
.B(net213),
.X(net219)
);

sky130_fd_sc_hd__a21o_2 c301(
.A1(in4),
.A2(net81),
.B1(net216),
.X(net220)
);

sky130_fd_sc_hd__mux4_1 c302(
.A0(net208),
.A1(net200),
.A2(out9),
.A3(net213),
.S0(net64),
.S1(net215),
.X(net221)
);

sky130_fd_sc_hd__or2b_1 c303(
.A(net219),
.B_N(net656),
.X(net222)
);

sky130_fd_sc_hd__mux4_2 c304(
.A0(net216),
.A1(net219),
.A2(net91),
.A3(net207),
.S0(net105),
.S1(net97),
.X(net223)
);

sky130_fd_sc_hd__buf_2 c305(
.A(net648),
.X(net224)
);

sky130_fd_sc_hd__mux4_1 c306(
.A0(net223),
.A1(net224),
.A2(net217),
.A3(in25),
.S0(net207),
.S1(net103),
.X(net225)
);

sky130_fd_sc_hd__o21ba_1 c307(
.A1(net224),
.A2(net216),
.B1_N(net219),
.X(net226)
);

sky130_fd_sc_hd__o21a_1 c308(
.A1(in14),
.A2(net102),
.B1(net190),
.X(net227)
);

sky130_fd_sc_hd__nand2b_2 c309(
.A_N(net92),
.B(net227),
.Y(net228)
);

sky130_fd_sc_hd__o21ba_4 c310(
.A1(net100),
.A2(net113),
.B1_N(in48),
.X(net229)
);

sky130_fd_sc_hd__or2b_1 c311(
.A(net207),
.B_N(out38),
.X(net230)
);

sky130_fd_sc_hd__nand2b_1 c312(
.A_N(in44),
.B(net210),
.Y(net231)
);

sky130_fd_sc_hd__nor2_4 c313(
.A(net227),
.B(in28),
.Y(net232)
);

sky130_fd_sc_hd__or2b_2 c314(
.A(net121),
.B_N(net194),
.X(net233)
);

sky130_fd_sc_hd__a21boi_2 c315(
.A1(net228),
.A2(net69),
.B1_N(net233),
.Y(net234)
);

sky130_fd_sc_hd__a311oi_4 c316(
.A1(net69),
.A2(net119),
.A3(in57),
.B1(net108),
.C1(net232),
.Y(net235)
);

sky130_fd_sc_hd__o21ai_0 c317(
.A1(net229),
.A2(net210),
.B1(net232),
.Y(net236)
);

sky130_fd_sc_hd__nor2b_1 c318(
.A(net190),
.B_N(net229),
.Y(out35)
);

sky130_fd_sc_hd__a21o_2 c319(
.A1(net235),
.A2(net193),
.B1(net234),
.X(net237)
);

sky130_fd_sc_hd__a311o_4 c320(
.A1(in28),
.A2(net233),
.A3(net210),
.B1(net230),
.C1(out35),
.X(net238)
);

sky130_fd_sc_hd__buf_8 c321(
.A(net639),
.X(net239)
);

sky130_fd_sc_hd__dfbbn_2 c322(
.D(net237),
.RESET_B(net235),
.SET_B(net233),
.CLK_N(clk),
.Q(net241),
.Q_N(net240)
);

sky130_fd_sc_hd__mux2_8 c323(
.A0(net231),
.A1(net234),
.S(net235),
.X(net242)
);

sky130_fd_sc_hd__a21bo_2 c324(
.A1(net238),
.A2(net231),
.B1_N(net219),
.X(net243)
);

sky130_fd_sc_hd__dfbbp_1 c325(
.D(net243),
.RESET_B(out35),
.SET_B(net230),
.CLK(clk),
.Q(out39),
.Q_N(net244)
);

sky130_fd_sc_hd__clkbuf_4 c326(
.A(net640),
.X(net245)
);

sky130_fd_sc_hd__a311oi_4 c327(
.A1(in57),
.A2(net125),
.A3(net113),
.B1(net234),
.C1(net90),
.Y(net246)
);

sky130_fd_sc_hd__sdfxbp_1 c328(
.D(net246),
.SCD(net231),
.SCE(net244),
.CLK(clk),
.Q(net248),
.Q_N(net247)
);

sky130_fd_sc_hd__sdfxbp_2 c329(
.D(net242),
.SCD(net245),
.SCE(out39),
.CLK(clk),
.Q(net250),
.Q_N(net249)
);

sky130_fd_sc_hd__nand2_4 c330(
.A(in47),
.B(in45),
.Y(net251)
);

sky130_fd_sc_hd__nand2b_1 c331(
.A_N(net145),
.B(net16),
.Y(net252)
);

sky130_fd_sc_hd__or2b_1 c332(
.A(in10),
.B_N(net16),
.X(net253)
);

sky130_fd_sc_hd__nor2b_1 c333(
.A(net251),
.B_N(net230),
.Y(net254)
);

sky130_fd_sc_hd__nor2_2 c334(
.A(net230),
.B(net249),
.Y(net255)
);

sky130_fd_sc_hd__inv_6 c335(
.A(net628),
.Y(net256)
);

sky130_fd_sc_hd__a211o_4 c336(
.A1(net142),
.A2(net255),
.B1(net134),
.C1(net234),
.X(net257)
);

sky130_fd_sc_hd__nand2b_2 c337(
.A_N(net150),
.B(net256),
.Y(net258)
);

sky130_fd_sc_hd__clkinv_2 c338(
.A(net627),
.Y(net259)
);

sky130_fd_sc_hd__and2_0 c339(
.A(net218),
.B(out25),
.X(out31)
);

sky130_fd_sc_hd__and2_0 c340(
.A(net256),
.B(net236),
.X(net260)
);

sky130_fd_sc_hd__or2b_1 c341(
.A(in48),
.B_N(out25),
.X(out61)
);

sky130_fd_sc_hd__clkbuf_16 c342(
.A(net650),
.X(net261)
);

sky130_fd_sc_hd__nand2b_4 c343(
.A_N(net261),
.B(net253),
.Y(out18)
);

sky130_fd_sc_hd__and2b_1 c344(
.A_N(net255),
.B(out61),
.X(net262)
);

sky130_fd_sc_hd__a21bo_4 c345(
.A1(net252),
.A2(out9),
.B1_N(net84),
.X(out29)
);

sky130_fd_sc_hd__nand2b_2 c346(
.A_N(net235),
.B(net253),
.Y(out37)
);

sky130_fd_sc_hd__nand2_2 c347(
.A(net260),
.B(net71),
.Y(net263)
);

sky130_fd_sc_hd__dfrtp_1 c348(
.D(net102),
.RESET_B(out37),
.CLK(clk),
.Q(net264)
);

sky130_fd_sc_hd__dfrtp_2 c349(
.D(net127),
.RESET_B(out37),
.CLK(clk),
.Q(net265)
);

sky130_fd_sc_hd__and2_2 c350(
.A(net119),
.B(net254),
.X(net266)
);

sky130_fd_sc_hd__mux4_2 c351(
.A0(net262),
.A1(net264),
.A2(net266),
.A3(out37),
.S0(net200),
.S1(net149),
.X(net267)
);

sky130_fd_sc_hd__a21bo_1 c352(
.A1(net259),
.A2(net240),
.B1_N(net159),
.X(out23)
);

sky130_fd_sc_hd__nor2b_1 c353(
.A(net103),
.B_N(out35),
.Y(net268)
);

sky130_fd_sc_hd__nor2b_2 c354(
.A(net40),
.B_N(net164),
.Y(net269)
);

sky130_fd_sc_hd__mux2_8 c355(
.A0(in27),
.A1(in26),
.S(out18),
.X(out52)
);

sky130_fd_sc_hd__nand2b_2 c356(
.A_N(net133),
.B(net97),
.Y(net270)
);

sky130_fd_sc_hd__sdfxtp_1 c357(
.D(net148),
.SCD(out22),
.SCE(net131),
.CLK(clk),
.Q(out56)
);

sky130_fd_sc_hd__and2b_4 c358(
.A_N(net166),
.B(net148),
.X(net271)
);

sky130_fd_sc_hd__sdfxtp_2 c359(
.D(net270),
.SCD(net131),
.SCE(in26),
.CLK(clk),
.Q(net272)
);

sky130_fd_sc_hd__inv_6 c360(
.A(net619),
.Y(net273)
);

sky130_fd_sc_hd__nand2_2 c361(
.A(net241),
.B(in27),
.Y(net274)
);

sky130_fd_sc_hd__buf_1 c362(
.A(net618),
.X(out26)
);

sky130_fd_sc_hd__or2_4 c363(
.A(net268),
.B(net30),
.X(net275)
);

sky130_fd_sc_hd__nor2b_2 c364(
.A(net274),
.B_N(net108),
.Y(net276)
);

sky130_fd_sc_hd__nand2b_2 c365(
.A_N(net33),
.B(net108),
.Y(net277)
);

sky130_fd_sc_hd__a21bo_1 c366(
.A1(net273),
.A2(net103),
.B1_N(net268),
.X(net278)
);

sky130_fd_sc_hd__and2b_2 c367(
.A_N(net277),
.B(net259),
.X(net279)
);

sky130_fd_sc_hd__a21boi_1 c368(
.A1(net276),
.A2(net271),
.B1_N(net84),
.Y(out50)
);

sky130_fd_sc_hd__mux4_4 c369(
.A0(net278),
.A1(net275),
.A2(net33),
.A3(out18),
.S0(net153),
.S1(out31),
.X(net280)
);

sky130_fd_sc_hd__sdfxtp_4 c370(
.D(net159),
.SCD(net280),
.SCE(in21),
.CLK(clk),
.Q(out55)
);

sky130_fd_sc_hd__and2_1 c371(
.A(net271),
.B(out35),
.X(net281)
);

sky130_fd_sc_hd__dfrtp_4 c372(
.D(net281),
.RESET_B(out39),
.CLK(clk),
.Q(net282)
);

sky130_fd_sc_hd__nand2_4 c373(
.A(net153),
.B(net282),
.Y(net283)
);

sky130_fd_sc_hd__mux4_4 c392(
.A0(net233),
.A1(net181),
.A2(out51),
.A3(out3),
.S0(out54),
.S1(out25),
.X(net284)
);

sky130_fd_sc_hd__mux4_4 c393(
.A0(net2),
.A1(out57),
.A2(out1),
.A3(net284),
.S0(out33),
.S1(out9),
.X(net285)
);

sky130_fd_sc_hd__mux4_1 c394(
.A0(net272),
.A1(out54),
.A2(out50),
.A3(out47),
.S0(out59),
.S1(out45),
.X(net286)
);

sky130_fd_sc_hd__mux4_2 c395(
.A0(net284),
.A1(in6),
.A2(out6),
.A3(net233),
.S0(out54),
.S1(out27),
.X(out60)
);

sky130_fd_sc_hd__nand2b_2 c396(
.A_N(net198),
.B(net74),
.Y(net287)
);

sky130_fd_sc_hd__inv_1 c397(
.A(net615),
.Y(net288)
);

sky130_fd_sc_hd__and2_4 c398(
.A(net202),
.B(net198),
.X(net289)
);

sky130_fd_sc_hd__nor2b_2 c399(
.A(net288),
.B_N(net188),
.Y(net290)
);

sky130_fd_sc_hd__or2b_1 c400(
.A(net201),
.B_N(net198),
.X(net291)
);

sky130_fd_sc_hd__and2_4 c401(
.A(in13),
.B(net291),
.X(net292)
);

sky130_fd_sc_hd__nand2_2 c402(
.A(in19),
.B(in0),
.Y(net293)
);

sky130_fd_sc_hd__and2b_2 c403(
.A_N(net290),
.B(net293),
.X(net294)
);

sky130_fd_sc_hd__buf_16 c404(
.A(net615),
.X(net295)
);

sky130_fd_sc_hd__nor2b_1 c405(
.A(net76),
.B_N(net295),
.Y(net296)
);

sky130_fd_sc_hd__clkinv_1 c406(
.A(net646),
.Y(net297)
);

sky130_fd_sc_hd__dfbbn_1 c407(
.D(net292),
.RESET_B(net294),
.SET_B(net295),
.CLK_N(clk),
.Q(net299),
.Q_N(net298)
);

sky130_fd_sc_hd__and2_2 c408(
.A(net74),
.B(net194),
.X(net300)
);

sky130_fd_sc_hd__mux4_1 c409(
.A0(net287),
.A1(net200),
.A2(net296),
.A3(net295),
.S0(net298),
.S1(net297),
.X(net301)
);

sky130_fd_sc_hd__mux2_8 c410(
.A0(net291),
.A1(net187),
.S(net295),
.X(net302)
);

sky130_fd_sc_hd__nor2_2 c411(
.A(net297),
.B(net295),
.Y(net303)
);

sky130_fd_sc_hd__a311o_1 c412(
.A1(net293),
.A2(net202),
.A3(net295),
.B1(net298),
.C1(net287),
.X(net304)
);

sky130_fd_sc_hd__dfsbp_1 c413(
.D(net300),
.SET_B(net205),
.CLK(clk),
.Q(net305)
);

sky130_fd_sc_hd__o21a_4 c414(
.A1(net305),
.A2(net295),
.B1(net303),
.X(net306)
);

sky130_fd_sc_hd__a21o_4 c415(
.A1(net295),
.A2(net296),
.B1(net198),
.X(net307)
);

sky130_fd_sc_hd__dfsbp_2 c416(
.D(net302),
.SET_B(net76),
.CLK(clk),
.Q(net309),
.Q_N(net308)
);

sky130_fd_sc_hd__dfbbn_2 c417(
.D(net296),
.RESET_B(net304),
.SET_B(net308),
.CLK_N(clk),
.Q(net311),
.Q_N(net310)
);

sky130_fd_sc_hd__buf_1 c418(
.A(net633),
.X(net312)
);

sky130_fd_sc_hd__or2b_4 c419(
.A(net94),
.B_N(net299),
.X(net313)
);

sky130_fd_sc_hd__nand2_1 c420(
.A(net211),
.B(net204),
.Y(net314)
);

sky130_fd_sc_hd__clkbuf_8 c421(
.A(net633),
.X(net315)
);

sky130_fd_sc_hd__or2_4 c422(
.A(net314),
.B(net203),
.X(net316)
);

sky130_fd_sc_hd__and2_2 c423(
.A(net316),
.B(net313),
.X(net317)
);

sky130_fd_sc_hd__inv_8 c424(
.A(net647),
.Y(net318)
);

sky130_fd_sc_hd__or2b_4 c425(
.A(net220),
.B_N(net315),
.X(net319)
);

sky130_fd_sc_hd__and2_4 c426(
.A(net296),
.B(net311),
.X(net320)
);

sky130_fd_sc_hd__nand2_2 c427(
.A(net313),
.B(net312),
.Y(net321)
);

sky130_fd_sc_hd__dfstp_1 c428(
.D(net319),
.SET_B(net320),
.CLK(clk),
.Q(net322)
);

sky130_fd_sc_hd__dfstp_2 c429(
.D(net315),
.SET_B(net319),
.CLK(clk),
.Q(net323)
);

sky130_fd_sc_hd__nand2_4 c430(
.A(net322),
.B(net94),
.Y(net324)
);

sky130_fd_sc_hd__dfstp_4 c431(
.D(net319),
.SET_B(net657),
.CLK(clk),
.Q(net325)
);

sky130_fd_sc_hd__nor2_2 c432(
.A(net321),
.B(net314),
.Y(out43)
);

sky130_fd_sc_hd__nor2_4 c433(
.A(net64),
.B(net322),
.Y(net326)
);

sky130_fd_sc_hd__nor2_1 c434(
.A(net325),
.B(net314),
.Y(net327)
);

sky130_fd_sc_hd__nand2b_1 c435(
.A_N(net312),
.B(net313),
.Y(net328)
);

sky130_fd_sc_hd__a21boi_1 c436(
.A1(net312),
.A2(net324),
.B1_N(net328),
.Y(net329)
);

sky130_fd_sc_hd__nor2b_2 c437(
.A(net327),
.B_N(net329),
.Y(net330)
);

sky130_fd_sc_hd__and2b_4 c438(
.A_N(net328),
.B(net220),
.X(net331)
);

sky130_fd_sc_hd__sdfbbp_1 c439(
.D(net91),
.RESET_B(net315),
.SCD(net331),
.SCE(net313),
.SET_B(out9),
.CLK(clk),
.Q(net332)
);

sky130_fd_sc_hd__sdfrbp_2 c440(
.D(net239),
.RESET_B(net331),
.SCD(net105),
.SCE(net294),
.CLK(clk),
.Q(net334),
.Q_N(net333)
);

sky130_fd_sc_hd__a211o_2 c441(
.A1(net324),
.A2(net334),
.B1(net93),
.C1(net236),
.X(net335)
);

sky130_fd_sc_hd__nor2b_1 c442(
.A(net228),
.B_N(net333),
.Y(net336)
);

sky130_fd_sc_hd__o21bai_1 c443(
.A1(net306),
.A2(net335),
.B1_N(net325),
.Y(net337)
);

sky130_fd_sc_hd__nand2b_1 c444(
.A_N(net194),
.B(net236),
.Y(net338)
);

sky130_fd_sc_hd__o21ba_1 c445(
.A1(net329),
.A2(net313),
.B1_N(net232),
.X(net339)
);

sky130_fd_sc_hd__clkbuf_4 c446(
.A(net638),
.X(net340)
);

sky130_fd_sc_hd__and2b_1 c447(
.A_N(net309),
.B(net306),
.X(net341)
);

sky130_fd_sc_hd__and2_1 c448(
.A(net227),
.B(net217),
.X(net342)
);

sky130_fd_sc_hd__a21boi_4 c449(
.A1(net232),
.A2(net247),
.B1_N(net323),
.Y(net343)
);

sky130_fd_sc_hd__o21ai_4 c450(
.A1(net124),
.A2(net342),
.B1(net336),
.Y(net344)
);

sky130_fd_sc_hd__a211oi_4 c451(
.A1(net338),
.A2(net108),
.B1(net294),
.C1(in25),
.Y(net345)
);

sky130_fd_sc_hd__and2_2 c452(
.A(net344),
.B(net341),
.X(net346)
);

sky130_fd_sc_hd__and2_1 c453(
.A(net248),
.B(net239),
.X(net347)
);

sky130_fd_sc_hd__and2b_4 c454(
.A_N(net105),
.B(net232),
.X(net348)
);

sky130_fd_sc_hd__inv_8 c455(
.A(net637),
.Y(net349)
);

sky130_fd_sc_hd__a211o_4 c456(
.A1(net347),
.A2(net344),
.B1(net348),
.C1(net227),
.X(net350)
);

sky130_fd_sc_hd__dfbbp_1 c457(
.D(net346),
.RESET_B(net349),
.SET_B(net350),
.CLK(clk),
.Q(net352),
.Q_N(net351)
);

sky130_fd_sc_hd__sdfrtn_1 c458(
.D(net345),
.RESET_B(net348),
.SCD(net93),
.SCE(in55),
.CLK_N(clk),
.Q(out17)
);

sky130_fd_sc_hd__mux4_4 c459(
.A0(net336),
.A1(net351),
.A2(net333),
.A3(net124),
.S0(net335),
.S1(net348),
.X(net353)
);

sky130_fd_sc_hd__mux4_4 c460(
.A0(net353),
.A1(net323),
.A2(net344),
.A3(net342),
.S0(net348),
.S1(net113),
.X(net354)
);

sky130_fd_sc_hd__or2_1 c461(
.A(net348),
.B(net352),
.X(net355)
);

sky130_fd_sc_hd__nor2_1 c462(
.A(net200),
.B(net196),
.Y(out8)
);

sky130_fd_sc_hd__sdfbbn_1 c463(
.D(net332),
.RESET_B(out37),
.SCD(in6),
.SCE(net236),
.SET_B(net16),
.CLK_N(clk),
.Q(net357),
.Q_N(net356)
);

sky130_fd_sc_hd__clkinv_16 c464(
.A(net623),
.Y(net358)
);

sky130_fd_sc_hd__or2_4 c465(
.A(net357),
.B(net658),
.X(net359)
);

sky130_fd_sc_hd__or2b_4 c466(
.A(net250),
.B_N(net657),
.X(net360)
);

sky130_fd_sc_hd__nor2b_1 c467(
.A(net357),
.B_N(net313),
.Y(net361)
);

sky130_fd_sc_hd__or2b_2 c468(
.A(net358),
.B_N(net357),
.X(net362)
);

sky130_fd_sc_hd__nand2_2 c469(
.A(net245),
.B(in55),
.Y(net363)
);

sky130_fd_sc_hd__a21boi_1 c470(
.A1(net18),
.A2(net362),
.B1_N(net134),
.Y(out0)
);

sky130_fd_sc_hd__sdfxbp_1 c471(
.D(net335),
.SCD(out12),
.SCE(net346),
.CLK(clk),
.Q(net364)
);

sky130_fd_sc_hd__mux4_4 c472(
.A0(net217),
.A1(net134),
.A2(out31),
.A3(in55),
.S0(net356),
.S1(net113),
.X(net365)
);

sky130_fd_sc_hd__mux4_4 c473(
.A0(net364),
.A1(net363),
.A2(net131),
.A3(net356),
.S0(net143),
.S1(net365),
.X(net366)
);

sky130_fd_sc_hd__nor2_2 c474(
.A(out25),
.B(net657),
.Y(net367)
);

sky130_fd_sc_hd__or2b_1 c475(
.A(net361),
.B_N(net135),
.X(net368)
);

sky130_fd_sc_hd__nand2b_1 c476(
.A_N(net236),
.B(net368),
.Y(net369)
);

sky130_fd_sc_hd__a211oi_1 c477(
.A1(net363),
.A2(in1),
.B1(net234),
.C1(net661),
.Y(net370)
);

sky130_fd_sc_hd__inv_16 c478(
.A(net624),
.Y(net371)
);

sky130_fd_sc_hd__sdfxbp_2 c479(
.D(net359),
.SCD(net370),
.SCE(net134),
.CLK(clk),
.Q(net373),
.Q_N(net372)
);

sky130_fd_sc_hd__mux2_2 c480(
.A0(net357),
.A1(net362),
.S(net661),
.X(out13)
);

sky130_fd_sc_hd__nand2_4 c481(
.A(net368),
.B(net306),
.Y(net374)
);

sky130_fd_sc_hd__mux4_4 c482(
.A0(net365),
.A1(net374),
.A2(net372),
.A3(net356),
.S0(net18),
.S1(net660),
.X(net375)
);

sky130_fd_sc_hd__mux4_1 c483(
.A0(net113),
.A1(net374),
.A2(net266),
.A3(net356),
.S0(net362),
.S1(net662),
.X(out21)
);

sky130_fd_sc_hd__or2_4 c484(
.A(net334),
.B(out38),
.X(net376)
);

sky130_fd_sc_hd__and2_0 c485(
.A(net339),
.B(net199),
.X(net377)
);

sky130_fd_sc_hd__nor2b_4 c486(
.A(net219),
.B_N(out11),
.Y(net378)
);

sky130_fd_sc_hd__a21boi_0 c487(
.A1(net108),
.A2(out29),
.B1_N(out16),
.Y(net379)
);

sky130_fd_sc_hd__sdfbbn_2 c488(
.D(net362),
.RESET_B(net199),
.SCD(net90),
.SCE(net378),
.SET_B(net341),
.CLK_N(clk),
.Q(net381),
.Q_N(net380)
);

sky130_fd_sc_hd__mux4_4 c489(
.A0(net371),
.A1(net164),
.A2(out35),
.A3(net378),
.S0(net244),
.S1(out16),
.X(net382)
);

sky130_fd_sc_hd__and2_4 c490(
.A(net376),
.B(net164),
.X(net383)
);

sky130_fd_sc_hd__o21ba_1 c491(
.A1(net144),
.A2(net135),
.B1_N(net32),
.X(net384)
);

sky130_fd_sc_hd__a211oi_4 c492(
.A1(net377),
.A2(out43),
.B1(in55),
.C1(out11),
.Y(net385)
);

sky130_fd_sc_hd__clkinv_2 c493(
.A(net634),
.Y(net386)
);

sky130_fd_sc_hd__buf_12 c494(
.A(net635),
.X(out41)
);

sky130_fd_sc_hd__sdfxtp_1 c495(
.D(net134),
.SCD(net383),
.SCE(net378),
.CLK(clk),
.Q(net387)
);

sky130_fd_sc_hd__mux4_1 c496(
.A0(net342),
.A1(net16),
.A2(out22),
.A3(net385),
.S0(out18),
.S1(net383),
.X(net388)
);

sky130_fd_sc_hd__sdfxtp_2 c497(
.D(net283),
.SCD(net377),
.SCE(net362),
.CLK(clk),
.Q(net389)
);

sky130_fd_sc_hd__a21boi_4 c498(
.A1(net135),
.A2(out31),
.B1_N(out30),
.Y(net390)
);

sky130_fd_sc_hd__or2_2 c499(
.A(in55),
.B(net663),
.X(net391)
);

sky130_fd_sc_hd__sdfxtp_4 c500(
.D(net390),
.SCD(net381),
.SCE(out25),
.CLK(clk),
.Q(net392)
);

sky130_fd_sc_hd__nand2b_2 c501(
.A_N(net16),
.B(net391),
.Y(net393)
);

sky130_fd_sc_hd__nor2_4 c502(
.A(net386),
.B(net393),
.Y(net394)
);

sky130_fd_sc_hd__a21bo_4 c503(
.A1(net384),
.A2(out18),
.B1_N(net326),
.X(net395)
);

sky130_fd_sc_hd__dfbbn_1 c504(
.D(net379),
.RESET_B(net392),
.SET_B(out26),
.CLK_N(clk),
.Q(net397),
.Q_N(net396)
);

sky130_fd_sc_hd__dfbbn_2 c505(
.D(net396),
.RESET_B(net385),
.SET_B(net664),
.CLK_N(clk),
.Q(net399),
.Q_N(net398)
);

sky130_fd_sc_hd__clkinv_1 c528(
.A(net645),
.Y(net400)
);

sky130_fd_sc_hd__and2b_2 c529(
.A_N(net293),
.B(net288),
.X(net401)
);

sky130_fd_sc_hd__nand2b_1 c530(
.A_N(net401),
.B(net310),
.Y(net402)
);

sky130_fd_sc_hd__or2_2 c531(
.A(net402),
.B(net400),
.X(net403)
);

sky130_fd_sc_hd__nand2_2 c532(
.A(in12),
.B(net401),
.Y(net404)
);

sky130_fd_sc_hd__clkinv_4 c533(
.A(net645),
.Y(net405)
);

sky130_fd_sc_hd__and2_1 c534(
.A(net402),
.B(net294),
.X(net406)
);

sky130_fd_sc_hd__nand2b_1 c535(
.A_N(net404),
.B(net303),
.Y(net407)
);

sky130_fd_sc_hd__and2_0 c536(
.A(net404),
.B(net291),
.X(net408)
);

sky130_fd_sc_hd__and2_1 c537(
.A(net303),
.B(net402),
.X(net409)
);

sky130_fd_sc_hd__or2b_4 c538(
.A(in0),
.B_N(net409),
.X(net410)
);

sky130_fd_sc_hd__nor2b_2 c539(
.A(net407),
.B_N(net188),
.Y(net411)
);

sky130_fd_sc_hd__nand2b_1 c540(
.A_N(net409),
.B(in12),
.Y(net412)
);

sky130_fd_sc_hd__nor2_4 c541(
.A(net406),
.B(net411),
.Y(net413)
);

sky130_fd_sc_hd__nor2b_4 c542(
.A(net410),
.B_N(net411),
.Y(net414)
);

sky130_fd_sc_hd__dfbbp_1 c543(
.D(net408),
.RESET_B(net410),
.SET_B(net404),
.CLK(clk),
.Q(net416),
.Q_N(net415)
);

sky130_fd_sc_hd__a21o_1 c544(
.A1(net412),
.A2(net411),
.B1(net188),
.X(net417)
);

sky130_fd_sc_hd__nand2b_4 c545(
.A_N(net288),
.B(net204),
.Y(net418)
);

sky130_fd_sc_hd__nand2b_2 c546(
.A_N(net413),
.B(net409),
.Y(net419)
);

sky130_fd_sc_hd__o21ai_1 c547(
.A1(net405),
.A2(net414),
.B1(net418),
.Y(net420)
);

sky130_fd_sc_hd__or2_4 c548(
.A(net414),
.B(net405),
.X(net421)
);

sky130_fd_sc_hd__a211o_4 c549(
.A1(net417),
.A2(net416),
.B1(net413),
.C1(net409),
.X(out19)
);

sky130_fd_sc_hd__o21ai_1 c550(
.A1(net208),
.A2(net188),
.B1(net294),
.Y(net422)
);

sky130_fd_sc_hd__dlygate4sd1_1 c551(
.A(net625),
.X(net423)
);

sky130_fd_sc_hd__and2b_4 c552(
.A_N(net409),
.B(net314),
.X(net424)
);

sky130_fd_sc_hd__a21o_1 c553(
.A1(net418),
.A2(net419),
.B1(net97),
.X(net425)
);

sky130_fd_sc_hd__and2b_2 c554(
.A_N(net406),
.B(net314),
.X(net426)
);

sky130_fd_sc_hd__nand2_2 c555(
.A(net416),
.B(net84),
.Y(net427)
);

sky130_fd_sc_hd__o21ai_1 c556(
.A1(net425),
.A2(net203),
.B1(out9),
.Y(net428)
);

sky130_fd_sc_hd__nor2_2 c557(
.A(net407),
.B(net107),
.Y(net429)
);

sky130_fd_sc_hd__o21a_4 c558(
.A1(net204),
.A2(net415),
.B1(net429),
.X(net430)
);

sky130_fd_sc_hd__sdfxbp_1 c559(
.D(net330),
.SCD(net425),
.SCE(net430),
.CLK(clk),
.Q(net432),
.Q_N(net431)
);

sky130_fd_sc_hd__mux2_4 c560(
.A0(net311),
.A1(in3),
.S(net211),
.X(net433)
);

sky130_fd_sc_hd__nand2b_1 c561(
.A_N(net423),
.B(net299),
.Y(net434)
);

sky130_fd_sc_hd__o21ba_2 c562(
.A1(net328),
.A2(net415),
.B1_N(net429),
.X(net435)
);

sky130_fd_sc_hd__mux2_2 c563(
.A0(net299),
.A1(net328),
.S(net433),
.X(net436)
);

sky130_fd_sc_hd__mux4_2 c564(
.A0(net424),
.A1(net434),
.A2(net431),
.A3(net429),
.S0(in12),
.S1(net436),
.X(net437)
);

sky130_fd_sc_hd__a21boi_2 c565(
.A1(net426),
.A2(net403),
.B1_N(net434),
.Y(net438)
);

sky130_fd_sc_hd__clkinv_2 c566(
.A(net626),
.Y(net439)
);

sky130_fd_sc_hd__sdfxbp_2 c567(
.D(net426),
.SCD(net193),
.SCE(net438),
.CLK(clk),
.Q(net441),
.Q_N(net440)
);

sky130_fd_sc_hd__sdfrtp_1 c568(
.D(net433),
.RESET_B(net435),
.SCD(net330),
.SCE(net419),
.CLK(clk),
.Q(net442)
);

sky130_fd_sc_hd__sdfxtp_1 c569(
.D(net434),
.SCD(net438),
.SCE(net441),
.CLK(clk),
.Q(net443)
);

sky130_fd_sc_hd__mux4_4 c570(
.A0(net400),
.A1(net318),
.A2(net439),
.A3(net420),
.S0(net314),
.S1(net440),
.X(out7)
);

sky130_fd_sc_hd__a211oi_4 c571(
.A1(net441),
.A2(net425),
.B1(net439),
.C1(net443),
.Y(net444)
);

sky130_fd_sc_hd__nand2_2 c572(
.A(net429),
.B(net344),
.Y(net445)
);

sky130_fd_sc_hd__inv_1 c573(
.A(net622),
.Y(net446)
);

sky130_fd_sc_hd__clkinv_16 c574(
.A(net622),
.Y(net447)
);

sky130_fd_sc_hd__mux4_1 c575(
.A0(in25),
.A1(net447),
.A2(net429),
.A3(in1),
.S0(net445),
.S1(net234),
.X(net448)
);

sky130_fd_sc_hd__and2_4 c576(
.A(net355),
.B(net665),
.X(net449)
);

sky130_fd_sc_hd__and2_0 c577(
.A(net442),
.B(net326),
.X(net450)
);

sky130_fd_sc_hd__nand2_1 c578(
.A(net450),
.B(net436),
.Y(net451)
);

sky130_fd_sc_hd__sdfxtp_2 c579(
.D(net446),
.SCD(net445),
.SCE(net438),
.CLK(clk),
.Q(net452)
);

sky130_fd_sc_hd__o21ai_0 c580(
.A1(net451),
.A2(net450),
.B1(net323),
.Y(net453)
);

sky130_fd_sc_hd__mux4_4 c581(
.A0(net453),
.A1(out19),
.A2(in55),
.A3(net427),
.S0(net450),
.S1(net413),
.X(net454)
);

sky130_fd_sc_hd__dlrbn_1 c582(
.D(net452),
.RESET_B(net445),
.GATE_N(clk),
.Q(net455)
);

sky130_fd_sc_hd__and2b_4 c583(
.A_N(net112),
.B(net323),
.X(net456)
);

sky130_fd_sc_hd__o21bai_2 c584(
.A1(net455),
.A2(net318),
.B1_N(net454),
.Y(net457)
);

sky130_fd_sc_hd__o21bai_1 c585(
.A1(net432),
.A2(net413),
.B1_N(net234),
.Y(net458)
);

sky130_fd_sc_hd__a21bo_2 c586(
.A1(net340),
.A2(net450),
.B1_N(net665),
.X(net459)
);

sky130_fd_sc_hd__dlrbn_2 c587(
.D(net458),
.RESET_B(net454),
.GATE_N(clk),
.Q(net460)
);

sky130_fd_sc_hd__a311o_4 c588(
.A1(net430),
.A2(net234),
.A3(net193),
.B1(net447),
.C1(in55),
.X(net461)
);

sky130_fd_sc_hd__dlrbp_1 c589(
.D(net457),
.RESET_B(net323),
.GATE(clk),
.Q(net463),
.Q_N(net462)
);

sky130_fd_sc_hd__sdfxtp_4 c590(
.D(net318),
.SCD(net461),
.SCE(net457),
.CLK(clk),
.Q(net464)
);

sky130_fd_sc_hd__a21o_1 c591(
.A1(net456),
.A2(net450),
.B1(out19),
.X(net465)
);

sky130_fd_sc_hd__or2_1 c592(
.A(net465),
.B(net460),
.X(net466)
);

sky130_fd_sc_hd__mux4_2 c593(
.A0(net323),
.A1(net454),
.A2(net462),
.A3(net464),
.S0(net442),
.S1(net466),
.X(net467)
);

sky130_fd_sc_hd__or2_1 c594(
.A(net436),
.B(out9),
.X(net468)
);

sky130_fd_sc_hd__inv_8 c595(
.A(net642),
.Y(net469)
);

sky130_fd_sc_hd__o21a_2 c596(
.A1(net373),
.A2(net447),
.B1(net97),
.X(net470)
);

sky130_fd_sc_hd__a211oi_1 c597(
.A1(net369),
.A2(net447),
.B1(out17),
.C1(net464),
.Y(net471)
);

sky130_fd_sc_hd__inv_1 c598(
.A(net643),
.Y(net472)
);

sky130_fd_sc_hd__o21a_2 c599(
.A1(net472),
.A2(net362),
.B1(out8),
.X(net473)
);

sky130_fd_sc_hd__a21oi_1 c600(
.A1(net473),
.A2(net469),
.B1(net326),
.Y(net474)
);

sky130_fd_sc_hd__o21bai_2 c601(
.A1(net464),
.A2(net468),
.B1_N(out9),
.Y(net475)
);

sky130_fd_sc_hd__dfbbn_1 c602(
.D(net474),
.RESET_B(in55),
.SET_B(net472),
.CLK_N(clk),
.Q(net476)
);

sky130_fd_sc_hd__dfbbn_2 c603(
.D(net289),
.RESET_B(net349),
.SET_B(net97),
.CLK_N(clk),
.Q(net477)
);

sky130_fd_sc_hd__a311o_4 c604(
.A1(net475),
.A2(net196),
.A3(net411),
.B1(net97),
.C1(net454),
.X(net478)
);

sky130_fd_sc_hd__a211oi_2 c605(
.A1(net470),
.A2(in1),
.B1(net472),
.C1(net411),
.Y(net479)
);

sky130_fd_sc_hd__and2_4 c606(
.A(net479),
.B(net454),
.X(net480)
);

sky130_fd_sc_hd__dfbbp_1 c607(
.D(net480),
.RESET_B(net475),
.SET_B(net466),
.CLK(clk),
.Q(out20),
.Q_N(net481)
);

sky130_fd_sc_hd__sdfxbp_1 c608(
.D(net471),
.SCD(net234),
.SCE(net436),
.CLK(clk),
.Q(net483),
.Q_N(net482)
);

sky130_fd_sc_hd__sdfbbp_1 c609(
.D(net437),
.RESET_B(out20),
.SCD(net480),
.SCE(net234),
.SET_B(out9),
.CLK(clk),
.Q(net485),
.Q_N(net484)
);

sky130_fd_sc_hd__sdfrtp_2 c610(
.D(net427),
.RESET_B(net474),
.SCD(net483),
.SCE(net472),
.CLK(clk),
.Q(net486)
);

sky130_fd_sc_hd__a311oi_4 c611(
.A1(net486),
.A2(net368),
.A3(net482),
.B1(net367),
.C1(out9),
.Y(net487)
);

sky130_fd_sc_hd__mux2_1 c612(
.A0(net477),
.A1(net71),
.S(net479),
.X(net488)
);

sky130_fd_sc_hd__mux4_2 c613(
.A0(net483),
.A1(net466),
.A2(net7),
.A3(net362),
.S0(net289),
.S1(net481),
.X(net489)
);

sky130_fd_sc_hd__sdfrtp_4 c614(
.D(net478),
.RESET_B(net487),
.SCD(net466),
.SCE(net454),
.CLK(clk),
.Q(out5)
);

sky130_fd_sc_hd__a21o_1 c615(
.A1(net468),
.A2(out5),
.B1(net411),
.X(net490)
);

sky130_fd_sc_hd__mux4_2 c616(
.A0(net131),
.A1(out13),
.A2(net30),
.A3(out16),
.S0(out9),
.S1(net84),
.X(net491)
);

sky130_fd_sc_hd__a211oi_1 c617(
.A1(net97),
.A2(net162),
.B1(net90),
.C1(net668),
.Y(net492)
);

sky130_fd_sc_hd__clkbuf_4 c618(
.A(net621),
.X(net493)
);

sky130_fd_sc_hd__a211oi_2 c619(
.A1(net397),
.A2(net459),
.B1(net97),
.C1(out11),
.Y(net494)
);

sky130_fd_sc_hd__a211o_4 c620(
.A1(net492),
.A2(net399),
.B1(out9),
.C1(net71),
.X(net495)
);

sky130_fd_sc_hd__a311o_4 c621(
.A1(net71),
.A2(net162),
.A3(net492),
.B1(net164),
.C1(net481),
.X(net496)
);

sky130_fd_sc_hd__o21ai_4 c622(
.A1(net30),
.A2(net279),
.B1(in11),
.Y(net497)
);

sky130_fd_sc_hd__inv_2 c623(
.A(net620),
.Y(out15)
);

sky130_fd_sc_hd__a21oi_2 c624(
.A1(net443),
.A2(net84),
.B1(out16),
.Y(net498)
);

sky130_fd_sc_hd__sdfxbp_2 c625(
.D(net387),
.SCD(net131),
.SCE(in11),
.CLK(clk),
.Q(net499)
);

sky130_fd_sc_hd__a311oi_2 c626(
.A1(net164),
.A2(net97),
.A3(net459),
.B1(net387),
.C1(net90),
.Y(net500)
);

sky130_fd_sc_hd__o21ai_2 c627(
.A1(net395),
.A2(net495),
.B1(net411),
.Y(net501)
);

sky130_fd_sc_hd__sdfsbp_1 c628(
.D(net498),
.SCD(net492),
.SCE(net443),
.SET_B(net341),
.CLK(clk),
.Q(out14)
);

sky130_fd_sc_hd__a311o_1 c629(
.A1(in6),
.A2(net398),
.A3(net326),
.B1(in17),
.C1(out12),
.X(net502)
);

sky130_fd_sc_hd__sdfxtp_1 c630(
.D(net499),
.SCD(net501),
.SCE(out0),
.CLK(clk),
.Q(net503)
);

sky130_fd_sc_hd__a21oi_1 c631(
.A1(net502),
.A2(net394),
.B1(net667),
.Y(out4)
);

sky130_fd_sc_hd__sdfsbp_2 c632(
.D(net494),
.SCD(net496),
.SCE(in1),
.SET_B(net503),
.CLK(clk),
.Q(net504)
);

sky130_fd_sc_hd__a21boi_1 c633(
.A1(in55),
.A2(net394),
.B1_N(net503),
.Y(net505)
);

sky130_fd_sc_hd__o21bai_4 c634(
.A1(net476),
.A2(net493),
.B1_N(out0),
.Y(net506)
);

sky130_fd_sc_hd__o21a_1 c635(
.A1(net301),
.A2(net506),
.B1(net495),
.X(net507)
);

sky130_fd_sc_hd__a211o_4 c636(
.A1(net411),
.A2(net90),
.B1(net506),
.C1(net164),
.X(out10)
);

sky130_fd_sc_hd__o21a_2 c637(
.A1(net503),
.A2(net505),
.B1(net504),
.X(net508)
);

sky130_fd_sc_hd__nand2b_2 c660(
.A_N(net291),
.B(in4),
.Y(net509)
);

sky130_fd_sc_hd__nor2_4 c661(
.A(net421),
.B(net420),
.Y(net510)
);

sky130_fd_sc_hd__clkbuf_4 c662(
.X(net511)
);

sky130_fd_sc_hd__or2b_4 c663(
.A(in2),
.B_N(in4),
.X(net512)
);

sky130_fd_sc_hd__clkinv_16 c664(
.A(net631),
.Y(net513)
);

sky130_fd_sc_hd__dlrbp_2 c665(
.D(in4),
.RESET_B(net292),
.GATE(clk),
.Q(net514)
);

sky130_fd_sc_hd__dlrtn_1 c666(
.D(net509),
.RESET_B(net188),
.GATE_N(clk),
.Q(net515)
);

sky130_fd_sc_hd__dlrtn_2 c667(
.D(net292),
.RESET_B(net421),
.GATE_N(clk),
.Q(net516)
);

sky130_fd_sc_hd__nand2b_4 c668(
.A_N(net516),
.B(net512),
.Y(net517)
);

sky130_fd_sc_hd__or2_2 c669(
.A(net513),
.B(net420),
.X(net518)
);

sky130_fd_sc_hd__dlrtn_4 c670(
.D(net518),
.RESET_B(net510),
.GATE_N(clk),
.Q(net519)
);

sky130_fd_sc_hd__or2b_4 c671(
.A(net519),
.B_N(net515),
.X(net520)
);

sky130_fd_sc_hd__a21bo_4 c672(
.A1(net517),
.A2(in4),
.B1_N(net519),
.X(net521)
);

sky130_fd_sc_hd__or2b_4 c673(
.A(net307),
.B_N(net403),
.X(net522)
);

sky130_fd_sc_hd__sdfxtp_2 c674(
.D(net187),
.SCD(net421),
.SCE(net510),
.CLK(clk),
.Q(net523)
);

sky130_fd_sc_hd__dlrtp_1 c675(
.D(net523),
.RESET_B(net510),
.GATE(clk),
.Q(net524)
);

sky130_fd_sc_hd__mux2_4 c676(
.A0(net524),
.A1(net511),
.S(net420),
.X(net525)
);

sky130_fd_sc_hd__a21bo_1 c677(
.A1(net514),
.A2(net522),
.B1_N(net524),
.X(net526)
);

sky130_fd_sc_hd__and2_2 c678(
.A(net521),
.B(net511),
.X(net527)
);

sky130_fd_sc_hd__nand2b_4 c679(
.A_N(net512),
.B(net527),
.Y(net528)
);

sky130_fd_sc_hd__sdfbbn_1 c680(
.D(net520),
.RESET_B(out19),
.SCD(net528),
.SCE(net527),
.SET_B(net525),
.CLK_N(clk),
.Q(net530),
.Q_N(net529)
);

sky130_fd_sc_hd__sdfbbn_2 c681(
.D(net526),
.RESET_B(net525),
.SCD(net527),
.SCE(net528),
.SET_B(net529),
.CLK_N(clk),
.Q(net532),
.Q_N(net531)
);

sky130_fd_sc_hd__nand2b_1 c682(
.A_N(net424),
.B(net528),
.Y(net533)
);

sky130_fd_sc_hd__sdfxtp_4 c683(
.D(net515),
.SCD(net444),
.SCE(net422),
.CLK(clk),
.Q(net534)
);

sky130_fd_sc_hd__o21bai_1 c684(
.A1(net527),
.A2(in6),
.B1_N(net424),
.Y(net535)
);

sky130_fd_sc_hd__clkbuf_16 c685(
.A(net641),
.X(net536)
);

sky130_fd_sc_hd__nor2b_4 c686(
.A(net188),
.B_N(net515),
.Y(net537)
);

sky130_fd_sc_hd__inv_12 c687(
.A(net641),
.Y(net538)
);

sky130_fd_sc_hd__and2b_2 c688(
.A_N(net420),
.B(net435),
.X(net539)
);

sky130_fd_sc_hd__dlrtp_2 c689(
.D(net534),
.RESET_B(net525),
.GATE(clk),
.Q(net540)
);

sky130_fd_sc_hd__dlrtp_4 c690(
.D(net535),
.RESET_B(net294),
.GATE(clk),
.Q(net541)
);

sky130_fd_sc_hd__nand2_1 c691(
.A(net403),
.B(net211),
.Y(net542)
);

sky130_fd_sc_hd__dfbbn_1 c692(
.D(net539),
.RESET_B(net542),
.SET_B(in4),
.CLK_N(clk),
.Q(net544),
.Q_N(net543)
);

sky130_fd_sc_hd__a21boi_0 c693(
.A1(net541),
.A2(net211),
.B1_N(net542),
.Y(net545)
);

sky130_fd_sc_hd__edfxbp_1 c694(
.D(net540),
.DE(net428),
.CLK(clk),
.Q(net546)
);

sky130_fd_sc_hd__edfxtp_1 c695(
.D(net546),
.DE(net525),
.CLK(clk),
.Q(net547)
);

sky130_fd_sc_hd__nand2_4 c696(
.A(net528),
.B(net542),
.Y(net548)
);

sky130_fd_sc_hd__sdfbbp_1 c697(
.D(net533),
.RESET_B(net534),
.SCD(net548),
.SCE(net527),
.SET_B(net536),
.CLK(clk),
.Q(net550),
.Q_N(net549)
);

sky130_fd_sc_hd__mux4_4 c698(
.A0(net203),
.A1(net294),
.A2(net548),
.A3(net534),
.S0(net549),
.S1(net527),
.X(net551)
);

sky130_fd_sc_hd__a21o_1 c699(
.A1(net548),
.A2(net551),
.B1(net542),
.X(net552)
);

sky130_fd_sc_hd__a311oi_1 c700(
.A1(net439),
.A2(net528),
.A3(net548),
.B1(net413),
.C1(net536),
.Y(net553)
);

sky130_fd_sc_hd__sdfbbn_1 c701(
.D(net428),
.RESET_B(net553),
.SCD(net548),
.SCE(net547),
.SET_B(net542),
.CLK_N(clk),
.Q(net555),
.Q_N(net554)
);

sky130_fd_sc_hd__sdfbbn_2 c702(
.D(net525),
.RESET_B(net552),
.SCD(net548),
.SCE(net551),
.SET_B(net534),
.CLK_N(clk),
.Q(net557),
.Q_N(net556)
);

sky130_fd_sc_hd__a311oi_1 c703(
.A1(net545),
.A2(net550),
.A3(net557),
.B1(net548),
.C1(net528),
.Y(net558)
);

sky130_fd_sc_hd__a21bo_2 c704(
.A1(net538),
.A2(net522),
.B1_N(net556),
.X(net559)
);

sky130_fd_sc_hd__nand2b_1 c705(
.A_N(net522),
.B(out19),
.Y(net560)
);

sky130_fd_sc_hd__a311o_4 c706(
.A1(net294),
.A2(net320),
.A3(net447),
.B1(net341),
.C1(net666),
.X(net561)
);

sky130_fd_sc_hd__dfbbn_2 c707(
.D(net337),
.RESET_B(net557),
.SET_B(net551),
.CLK_N(clk),
.Q(net562)
);

sky130_fd_sc_hd__buf_8 c708(
.A(net644),
.X(net563)
);

sky130_fd_sc_hd__a21bo_1 c709(
.A1(net320),
.A2(net559),
.B1_N(net529),
.X(net564)
);

sky130_fd_sc_hd__dfbbp_1 c710(
.D(net563),
.RESET_B(net564),
.SET_B(net659),
.CLK(clk),
.Q(net565)
);

sky130_fd_sc_hd__a21bo_2 c711(
.A1(net551),
.A2(net554),
.B1_N(net320),
.X(net566)
);

sky130_fd_sc_hd__sdfxbp_1 c712(
.D(net557),
.SCD(net564),
.SCE(net538),
.CLK(clk),
.Q(net567)
);

sky130_fd_sc_hd__nor2b_2 c713(
.A(in21),
.B_N(net565),
.Y(net568)
);

sky130_fd_sc_hd__sdfxbp_2 c714(
.D(net93),
.SCD(net517),
.SCE(net449),
.CLK(clk),
.Q(net569)
);

sky130_fd_sc_hd__a21o_2 c715(
.A1(net193),
.A2(net562),
.B1(net556),
.X(net570)
);

sky130_fd_sc_hd__sdfxtp_1 c716(
.D(net537),
.SCD(net532),
.SCE(net564),
.CLK(clk),
.Q(net571)
);

sky130_fd_sc_hd__clkbuf_2 c717(
.A(net644),
.X(net572)
);

sky130_fd_sc_hd__nor2b_4 c718(
.A(net435),
.B_N(net571),
.Y(net573)
);

sky130_fd_sc_hd__o21ai_2 c719(
.A1(net569),
.A2(net542),
.B1(net572),
.Y(net574)
);

sky130_fd_sc_hd__mux4_2 c720(
.A0(net560),
.A1(net574),
.A2(net517),
.A3(out19),
.S0(net564),
.S1(net572),
.X(net575)
);

sky130_fd_sc_hd__or2_1 c721(
.A(net542),
.B(net572),
.X(net576)
);

sky130_fd_sc_hd__o21ai_4 c722(
.A1(net555),
.A2(net572),
.B1(net669),
.Y(net577)
);

sky130_fd_sc_hd__sdlclkp_1 c723(
.GATE(net564),
.SCE(net566),
.CLK(clk),
.GCLK(net578)
);

sky130_fd_sc_hd__o21bai_4 c724(
.A1(net573),
.A2(net561),
.B1_N(net578),
.Y(net579)
);

sky130_fd_sc_hd__sdfxtp_2 c725(
.D(net570),
.SCD(net579),
.SCE(net435),
.CLK(clk),
.Q(net580)
);

sky130_fd_sc_hd__inv_4 c726(
.A(net614),
.Y(net581)
);

sky130_fd_sc_hd__clkinv_4 c727(
.A(net613),
.Y(net582)
);

sky130_fd_sc_hd__o21ai_4 c728(
.A1(net367),
.A2(net582),
.B1(out19),
.Y(net583)
);

sky130_fd_sc_hd__a21oi_4 c729(
.A1(net580),
.A2(net341),
.B1(net582),
.Y(net584)
);

sky130_fd_sc_hd__a21o_2 c730(
.A1(net547),
.A2(net572),
.B1(net7),
.X(net585)
);

sky130_fd_sc_hd__a311o_1 c731(
.A1(net582),
.A2(in6),
.A3(net196),
.B1(net536),
.C1(net7),
.X(net586)
);

sky130_fd_sc_hd__o21bai_4 c732(
.A1(net447),
.A2(net586),
.B1_N(net582),
.Y(net587)
);

sky130_fd_sc_hd__nand2b_4 c733(
.A_N(net536),
.B(net572),
.Y(net588)
);

sky130_fd_sc_hd__or2b_1 c734(
.A(net587),
.B_N(net7),
.X(net589)
);

sky130_fd_sc_hd__o21ba_4 c735(
.A1(net567),
.A2(net585),
.B1_N(net530),
.X(net590)
);

sky130_fd_sc_hd__o21bai_2 c736(
.A1(net583),
.A2(net582),
.B1_N(net484),
.Y(net591)
);

sky130_fd_sc_hd__sdfxtp_4 c737(
.D(net591),
.SCD(net590),
.SCE(net341),
.CLK(clk),
.Q(net592)
);

sky130_fd_sc_hd__mux4_2 c738(
.A0(net577),
.A1(net581),
.A2(net580),
.A3(net341),
.S0(net582),
.S1(in11),
.X(net593)
);

sky130_fd_sc_hd__a21o_1 c739(
.A1(net584),
.A2(net592),
.B1(net582),
.X(net594)
);

sky130_fd_sc_hd__a21o_1 c740(
.A1(net576),
.A2(net490),
.B1(net666),
.X(net595)
);

sky130_fd_sc_hd__o21ba_4 c741(
.A1(net254),
.A2(net594),
.B1_N(net582),
.X(net596)
);

sky130_fd_sc_hd__mux4_2 c742(
.A0(net532),
.A1(net588),
.A2(net447),
.A3(net582),
.S0(net572),
.S1(net7),
.X(net597)
);

sky130_fd_sc_hd__mux4_4 c743(
.A0(net264),
.A1(net490),
.A2(net597),
.A3(in11),
.S0(net580),
.S1(net591),
.X(net598)
);

sky130_fd_sc_hd__o21ba_1 c744(
.A1(net568),
.A2(net596),
.B1_N(net580),
.X(net599)
);

sky130_fd_sc_hd__dfbbn_1 c745(
.D(net589),
.RESET_B(net463),
.SET_B(net595),
.CLK_N(clk),
.Q(net600)
);

sky130_fd_sc_hd__o21a_1 c746(
.A1(net593),
.A2(net599),
.B1(net670),
.X(net601)
);

sky130_fd_sc_hd__o21bai_1 c747(
.A1(net601),
.A2(net597),
.B1_N(net7),
.Y(net602)
);

sky130_fd_sc_hd__a311oi_1 c748(
.A1(net196),
.A2(net544),
.A3(net459),
.B1(net602),
.C1(net341),
.Y(net603)
);

sky130_fd_sc_hd__a211o_2 c749(
.A1(net389),
.A2(net530),
.B1(net558),
.C1(net349),
.X(net604)
);

sky130_fd_sc_hd__sdfstp_1 c750(
.D(net485),
.SCD(net500),
.SCE(net530),
.SET_B(net459),
.CLK(clk),
.Q(net605)
);

sky130_fd_sc_hd__a311o_4 c751(
.A1(net341),
.A2(net603),
.A3(net605),
.B1(net459),
.C1(net389),
.X(net606)
);

sky130_fd_sc_hd__a211oi_4 c752(
.A1(net459),
.A2(net349),
.B1(net602),
.C1(net389),
.Y(net607)
);

sky130_fd_sc_hd__a311o_2 c753(
.A1(net607),
.A2(net605),
.A3(net508),
.B1(out19),
.C1(net389),
.X(net608)
);

sky130_fd_sc_hd__sdfbbp_1 c754(
.D(net606),
.RESET_B(net608),
.SCD(net459),
.SCE(net558),
.SET_B(net508),
.CLK(clk),
.Q(net609)
);

sky130_fd_sc_hd__sdfbbn_1 c755(
.D(net326),
.RESET_B(net609),
.SCD(net507),
.SCE(net389),
.SET_B(net608),
.CLK_N(clk),
.Q(net610)
);

sky130_fd_sc_hd__a311o_4 c756(
.A1(net604),
.A2(net610),
.A3(net600),
.B1(net341),
.C1(net543)
);

sky130_fd_sc_hd__dfbbn_2 merge757(
.D(net141),
.RESET_B(net134),
.SET_B(in7),
.CLK_N(clk),
.Q(net612),
.Q_N(net611)
);

sky130_fd_sc_hd__sdfbbn_2 merge758(
.D(net469),
.RESET_B(net346),
.SCD(net529),
.SCE(net488),
.SET_B(net531),
.CLK_N(clk),
.Q(net614),
.Q_N(net613)
);

sky130_fd_sc_hd__sdfstp_2 merge759(
.D(net205),
.SCD(out38),
.SCE(net292),
.SET_B(net290),
.CLK(clk),
.Q(net615)
);

sky130_fd_sc_hd__dfbbp_1 merge760(
.D(net129),
.RESET_B(net131),
.SET_B(in52),
.CLK(clk),
.Q(net617),
.Q_N(net616)
);

sky130_fd_sc_hd__sdfxbp_1 merge761(
.D(net269),
.SCD(out46),
.SCE(net265),
.CLK(clk),
.Q(net619),
.Q_N(net618)
);

sky130_fd_sc_hd__sdfbbp_1 merge762(
.D(net32),
.RESET_B(net378),
.SCD(out13),
.SCE(net497),
.SET_B(net482),
.CLK(clk),
.Q(net621),
.Q_N(net620)
);

sky130_fd_sc_hd__sdfstp_4 merge763(
.D(net445),
.SCD(net289),
.SCE(net65),
.SET_B(net350),
.CLK(clk),
.Q(net622)
);

sky130_fd_sc_hd__sdfbbn_1 merge764(
.D(net360),
.RESET_B(net365),
.SCD(net263),
.SCE(net349),
.SET_B(net342),
.CLK_N(clk),
.Q(net624),
.Q_N(net623)
);

sky130_fd_sc_hd__sdfbbn_2 merge765(
.D(net408),
.RESET_B(net438),
.SCD(net419),
.SCE(in17),
.SET_B(net330),
.CLK_N(clk),
.Q(net626),
.Q_N(net625)
);

sky130_fd_sc_hd__sedfxbp_1 merge766(
.D(net149),
.DE(net238),
.SCD(net257),
.SCE(net113),
.CLK(clk),
.Q(net628),
.Q_N(net627)
);

sky130_fd_sc_hd__sedfxbp_2 merge767(
.D(net52),
.DE(net172),
.SCD(net180),
.SCE(out42),
.CLK(clk),
.Q(net630),
.Q_N(net629)
);

sky130_fd_sc_hd__sdfxbp_2 merge768(
.D(net510),
.SCD(net413),
.Q(net511),
.CLK(clk),
.Q_N(net631)
);

sky130_fd_sc_hd__sdfxtp_1 merge769(
.D(net215),
.SCD(net200),
.SCE(net290),
.CLK(clk),
.Q(net633)
);

sky130_fd_sc_hd__sdfbbp_1 merge770(
.D(net380),
.RESET_B(out1),
.SCD(net385),
.SCE(net71),
.SET_B(net301),
.CLK(clk),
.Q(net635),
.Q_N(net634)
);

sky130_fd_sc_hd__sedfxtp_1 merge771(
.D(net14),
.DE(net43),
.SCD(net50),
.SCE(net53),
.CLK(clk),
.Q(net636)
);

sky130_fd_sc_hd__sdfbbn_1 merge772(
.D(net331),
.RESET_B(in21),
.SCD(in25),
.SCE(net343),
.SET_B(in3),
.CLK_N(clk),
.Q(net638),
.Q_N(net637)
);

sky130_fd_sc_hd__sdfbbn_2 merge773(
.D(net234),
.RESET_B(net237),
.SCD(net226),
.SCE(net236),
.SET_B(out35),
.CLK_N(clk),
.Q(net640),
.Q_N(net639)
);

sky130_fd_sc_hd__sedfxtp_2 merge774(
.D(net444),
.DE(net326),
.SCD(net422),
.SCE(net525),
.CLK(clk),
.Q(net641)
);

sky130_fd_sc_hd__sdfbbp_1 merge775(
.D(net266),
.RESET_B(out21),
.SCD(net438),
.SCE(net234),
.SET_B(net443),
.CLK(clk),
.Q(net643),
.Q_N(net642)
);

sky130_fd_sc_hd__sedfxtp_4 merge776(
.D(net461),
.DE(net413),
.SCD(net449),
.SCE(net564),
.CLK(clk),
.Q(net644)
);

sky130_fd_sc_hd__sdfxtp_2 merge777(
.D(net304),
.SCD(in0),
.SCE(net66),
.CLK(clk),
.Q(net645)
);

sky130_fd_sc_hd__sdfrbp_1 merge778(
.D(net317),
.RESET_B(net204),
.SCD(net289),
.SCE(net64),
.CLK(clk),
.Q(net647),
.Q_N(net646)
);

sky130_fd_sc_hd__sdfrbp_2 merge779(
.D(net205),
.RESET_B(net200),
.SCD(net222),
.SCE(net217),
.CLK(clk),
.Q(net649),
.Q_N(net648)
);

sky130_fd_sc_hd__sdfrtn_1 merge780(
.D(net258),
.RESET_B(net103),
.SCD(net140),
.SCE(net141),
.CLK_N(clk),
.Q(net650)
);

sky130_fd_sc_hd__sdfrtp_1 merge781(
.D(net139),
.RESET_B(net131),
.SCD(net9),
.SCE(net141),
.CLK(clk),
.Q(net651)
);

sky130_fd_sc_hd__dfxbp_1 s782(
.D(net44),
.CLK(clk),
.Q(out30),
.Q_N(net652)
);

sky130_fd_sc_hd__dfxbp_2 s783(
.D(net60),
.CLK(clk),
.Q(net654),
.Q_N(net653)
);

sky130_fd_sc_hd__dfxtp_1 s784(
.D(net168),
.CLK(clk),
.Q(net655)
);

sky130_fd_sc_hd__dfxtp_2 s785(
.D(net221),
.CLK(clk),
.Q(net656)
);

sky130_fd_sc_hd__dfxtp_4 s786(
.D(net225),
.CLK(clk),
.Q(net657)
);

sky130_fd_sc_hd__dlclkp_1 s787(
.GATE(net267),
.CLK(clk),
.GCLK(net658)
);

sky130_fd_sc_hd__dlclkp_2 s788(
.GATE(net285),
.CLK(clk),
.GCLK(out45)
);

sky130_fd_sc_hd__dlclkp_4 s789(
.GATE(net286),
.CLK(clk),
.GCLK(out27)
);

sky130_fd_sc_hd__dlxbn_1 s790(
.D(net354),
.GATE_N(clk),
.Q(net659)
);

sky130_fd_sc_hd__dlxbn_2 s791(
.D(net366),
.GATE_N(clk),
.Q(net661),
.Q_N(net660)
);

sky130_fd_sc_hd__dlxbp_1 s792(
.D(net375),
.GATE(clk),
.Q(net662)
);

sky130_fd_sc_hd__dlxtn_1 s793(
.D(net382),
.GATE_N(clk),
.Q(net663)
);

sky130_fd_sc_hd__dlxtn_2 s794(
.D(net388),
.GATE_N(clk),
.Q(net664)
);

sky130_fd_sc_hd__dlxtn_4 s795(
.D(net448),
.GATE_N(clk),
.Q(net665)
);

sky130_fd_sc_hd__dlxtp_1 s796(
.D(net467),
.GATE(clk),
.Q(net666)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s797(
.D(net489),
.SLEEP_B(clk),
.Q(net667)
);

sky130_fd_sc_hd__dfxbp_1 s798(
.D(net491),
.CLK(clk),
.Q(net668)
);

sky130_fd_sc_hd__dfxbp_2 s799(
.D(net575),
.CLK(clk),
.Q(net669)
);

sky130_fd_sc_hd__dfxtp_1 s800(
.D(net598),
.CLK(clk),
.Q(net670)
);


endmodule
