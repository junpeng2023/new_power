module netlist_0 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input in52,
	input in53,
	input in54,
	input in55,
	input in56,
	input in57,
	input in58,
	input in59,
	input in60,
	input in61,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51,
	output out52,
	output out53,
	output out54,
	output out55,
	output out56,
	output out57,
	output out58,
	output out59,
	output out60,
	output out61
);


wire clk;
wire net860;
wire net857;
wire net854;
wire net853;
wire net851;
wire net850;
wire net849;
wire net848;
wire net846;
wire net844;
wire net842;
wire net841;
wire out3;
wire net837;
wire out19;
wire net834;
wire net833;
wire net832;
wire net831;
wire net829;
wire net827;
wire net825;
wire net843;
wire net823;
wire net822;
wire net821;
wire net820;
wire net819;
wire net818;
wire net817;
wire net816;
wire net815;
wire out13;
wire net814;
wire net813;
wire net812;
wire net811;
wire net810;
wire net807;
wire out24;
wire net805;
wire net804;
wire net802;
wire net801;
wire net800;
wire net795;
wire net793;
wire net792;
wire out56;
wire net791;
wire net789;
wire net787;
wire net786;
wire net785;
wire net784;
wire net808;
wire net781;
wire net780;
wire out1;
wire net777;
wire net776;
wire net775;
wire net774;
wire out43;
wire net773;
wire net772;
wire net771;
wire net770;
wire net769;
wire net766;
wire out15;
wire net765;
wire net764;
wire net763;
wire net762;
wire out52;
wire net759;
wire net755;
wire net754;
wire net753;
wire out42;
wire net752;
wire net751;
wire out49;
wire net750;
wire net748;
wire net790;
wire net747;
wire net745;
wire net744;
wire net743;
wire net741;
wire net740;
wire net739;
wire net738;
wire net735;
wire net732;
wire net731;
wire net730;
wire net729;
wire net728;
wire net726;
wire net725;
wire net724;
wire net722;
wire net720;
wire net719;
wire net717;
wire net716;
wire net715;
wire net714;
wire net712;
wire net711;
wire net708;
wire net706;
wire net705;
wire out30;
wire net704;
wire net703;
wire net701;
wire net699;
wire out40;
wire net692;
wire net690;
wire net299;
wire net688;
wire net686;
wire net684;
wire net683;
wire out57;
wire net503;
wire net679;
wire net671;
wire net669;
wire net668;
wire net370;
wire net667;
wire net664;
wire net694;
wire net659;
wire out54;
wire in6;
wire net656;
wire net652;
wire net622;
wire net651;
wire net304;
wire net645;
wire net641;
wire net637;
wire net632;
wire net665;
wire net631;
wire net629;
wire net74;
wire net628;
wire net3;
wire net627;
wire net447;
wire net626;
wire net624;
wire net506;
wire net623;
wire net620;
wire in49;
wire net619;
wire net798;
wire net46;
wire net615;
wire net100;
wire net347;
wire net288;
wire net614;
wire net165;
wire net613;
wire net20;
wire net612;
wire net638;
wire net428;
wire net610;
wire out25;
wire net608;
wire net1;
wire net424;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire net782;
wire net601;
wire net596;
wire net384;
wire net482;
wire net595;
wire net592;
wire net588;
wire net587;
wire in4;
wire net583;
wire net707;
wire net582;
wire net158;
wire net584;
wire net581;
wire net336;
wire net579;
wire net577;
wire net576;
wire net209;
wire net569;
wire in41;
wire net567;
wire net696;
wire net794;
wire in30;
wire net566;
wire net565;
wire net39;
wire net562;
wire net559;
wire net556;
wire net647;
wire net555;
wire net159;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire in55;
wire net550;
wire net710;
wire net544;
wire net539;
wire net534;
wire net532;
wire net271;
wire net530;
wire net617;
wire net306;
wire net537;
wire net369;
wire net528;
wire net525;
wire net523;
wire net520;
wire net519;
wire out6;
wire out20;
wire net516;
wire net672;
wire net514;
wire net78;
wire net508;
wire net721;
wire net504;
wire net224;
wire net573;
wire net499;
wire net674;
wire net496;
wire net495;
wire net494;
wire net179;
wire in39;
wire net453;
wire net493;
wire net788;
wire net472;
wire net492;
wire net479;
wire net491;
wire net295;
wire net490;
wire net489;
wire net856;
wire net487;
wire net486;
wire net478;
wire net474;
wire net473;
wire net468;
wire net540;
wire net202;
wire net465;
wire out7;
wire net462;
wire net469;
wire net471;
wire net461;
wire net546;
wire net749;
wire net460;
wire out17;
wire net454;
wire net44;
wire net117;
wire net689;
wire net859;
wire net858;
wire net648;
wire net452;
wire net449;
wire net448;
wire net835;
wire out11;
wire net498;
wire net700;
wire net446;
wire net680;
wire net88;
wire net691;
wire net444;
wire in59;
wire net110;
wire net442;
wire net441;
wire net609;
wire net440;
wire net128;
wire net439;
wire out21;
wire net147;
wire net438;
wire net797;
wire net433;
wire net432;
wire out41;
wire net419;
wire net431;
wire net430;
wire net618;
wire net429;
wire net427;
wire net809;
wire net426;
wire net673;
wire net425;
wire net570;
wire out2;
wire net423;
wire net183;
wire net531;
wire net421;
wire net52;
wire net170;
wire net420;
wire net450;
wire net418;
wire net416;
wire net779;
wire net698;
wire net839;
wire out23;
wire net512;
wire net18;
wire out34;
wire net415;
wire net414;
wire net276;
wire net413;
wire net330;
wire net252;
wire net412;
wire net411;
wire net826;
wire net517;
wire net677;
wire net410;
wire net409;
wire net475;
wire net408;
wire net685;
wire net407;
wire net406;
wire net662;
wire net405;
wire net836;
wire net607;
wire net526;
wire net404;
wire net29;
wire net403;
wire net383;
wire net663;
wire net402;
wire net106;
wire net572;
wire net401;
wire net847;
wire net399;
wire net398;
wire net476;
wire net855;
wire net396;
wire net172;
wire net395;
wire net391;
wire net693;
wire net443;
wire net557;
wire net345;
wire net527;
wire net488;
wire net390;
wire out5;
wire net646;
wire net389;
wire net513;
wire net501;
wire out14;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net184;
wire net131;
wire net380;
wire net379;
wire net260;
wire net616;
wire net378;
wire net543;
wire net38;
wire net377;
wire net376;
wire net625;
wire net373;
wire net598;
wire net374;
wire net676;
wire net372;
wire net371;
wire net368;
wire net367;
wire net366;
wire net365;
wire net364;
wire net363;
wire net360;
wire out18;
wire net397;
wire net357;
wire net356;
wire net510;
wire net355;
wire net590;
wire net507;
wire net351;
wire net746;
wire net350;
wire net547;
wire net511;
wire net451;
wire net13;
wire net343;
wire net89;
wire net666;
wire net340;
wire net339;
wire net337;
wire net458;
wire net538;
wire net244;
wire net334;
wire net333;
wire net332;
wire net331;
wire net328;
wire net327;
wire net119;
wire net325;
wire net324;
wire net321;
wire net535;
wire net320;
wire net542;
wire net139;
wire net318;
wire out9;
wire net335;
wire net315;
wire net505;
wire net199;
wire out27;
wire net294;
wire net319;
wire net312;
wire net636;
wire net518;
wire in37;
wire net311;
wire net309;
wire net742;
wire net308;
wire net417;
wire out8;
wire net302;
wire net298;
wire net296;
wire in24;
wire net358;
wire net127;
wire net180;
wire net310;
wire net697;
wire net293;
wire net305;
wire net292;
wire net521;
wire net353;
wire net500;
wire net445;
wire net230;
wire out22;
wire net303;
wire net291;
wire net201;
wire net422;
wire net289;
wire in25;
wire net589;
wire net278;
wire net761;
wire net274;
wire net643;
wire net273;
wire net272;
wire net114;
wire net270;
wire in17;
wire net267;
wire net644;
wire net266;
wire net459;
wire net463;
wire net0;
wire net297;
wire net280;
wire net102;
wire net799;
wire net151;
wire net275;
wire net264;
wire net657;
wire net591;
wire net196;
wire net262;
wire net217;
wire net261;
wire net21;
wire net257;
wire net62;
wire net109;
wire net254;
wire net203;
wire net253;
wire net188;
wire net207;
wire out16;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire net767;
wire net111;
wire net124;
wire net242;
wire in26;
wire net661;
wire net194;
wire net241;
wire out38;
wire in29;
wire net240;
wire net238;
wire net286;
wire net153;
wire out61;
wire out10;
wire net142;
wire net234;
wire net232;
wire out12;
wire net226;
wire out32;
wire net568;
wire net375;
wire net223;
wire net524;
wire net575;
wire net382;
wire net852;
wire net548;
wire net259;
wire net222;
wire net31;
wire net219;
wire net578;
wire net210;
wire net326;
wire net213;
wire net208;
wire net649;
wire net205;
wire net678;
wire net633;
wire net122;
wire net197;
wire net840;
wire net483;
wire net193;
wire net192;
wire net737;
wire net190;
wire net630;
wire in20;
wire net189;
wire net246;
wire net783;
wire net186;
wire net152;
wire net126;
wire net113;
wire net284;
wire net655;
wire net563;
wire net464;
wire net549;
wire net182;
wire net258;
wire net176;
wire net342;
wire net17;
wire net437;
wire out44;
wire net580;
wire net133;
wire net175;
wire net80;
wire net173;
wire net195;
wire net41;
wire net104;
wire net8;
wire net381;
wire net218;
wire net300;
wire net169;
wire out58;
wire net828;
wire net485;
wire net344;
wire net168;
wire net167;
wire net509;
wire net58;
wire net221;
wire net166;
wire net269;
wire net97;
wire net434;
wire net204;
wire net200;
wire net621;
wire net162;
wire out60;
wire net497;
wire out45;
wire net161;
wire net285;
wire net160;
wire net316;
wire out31;
wire net150;
wire net149;
wire net695;
wire net148;
wire net178;
wire net239;
wire net144;
wire net322;
wire net758;
wire net143;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net806;
wire net561;
wire out29;
wire net137;
wire net136;
wire net456;
wire net135;
wire net255;
wire net157;
wire net177;
wire net349;
wire out51;
wire out48;
wire net134;
wire net250;
wire net225;
wire net132;
wire net130;
wire in12;
wire net103;
wire net481;
wire net120;
wire net392;
wire out0;
wire net164;
wire net687;
wire net642;
wire net268;
wire in7;
wire net756;
wire net400;
wire net82;
wire net2;
wire net123;
wire net282;
wire net71;
wire net229;
wire in43;
wire net108;
wire net107;
wire net99;
wire net6;
wire net457;
wire out50;
wire net348;
wire net341;
wire in52;
wire net96;
wire net466;
wire net118;
wire net94;
wire net90;
wire net803;
wire net174;
wire net277;
wire net639;
wire net81;
wire net75;
wire net231;
wire net329;
wire net212;
wire net653;
wire in5;
wire net14;
wire net77;
wire net600;
wire net236;
wire net76;
wire in42;
wire net354;
wire in38;
wire net736;
wire net198;
wire net467;
wire net101;
wire net9;
wire net571;
wire net73;
wire net60;
wire net564;
wire net154;
wire net84;
wire net237;
wire net682;
wire in46;
wire net85;
wire net72;
wire net116;
wire net69;
wire net67;
wire net98;
wire net522;
wire net436;
wire net541;
wire net323;
wire net15;
wire net279;
wire net64;
wire net63;
wire net681;
wire net61;
wire net59;
wire net248;
wire net477;
wire net156;
wire in10;
wire net228;
wire net675;
wire net56;
wire out53;
wire net55;
wire net214;
wire net53;
wire in48;
wire net660;
wire net838;
wire net359;
wire out28;
wire net640;
wire net50;
wire in31;
wire net129;
wire net65;
wire net597;
wire out55;
wire net185;
wire net155;
wire net338;
wire net599;
wire net112;
wire net650;
wire net79;
wire net585;
wire net560;
wire net45;
wire net502;
wire net235;
wire net830;
wire net49;
wire out39;
wire net594;
wire in50;
wire net215;
wire net484;
wire in8;
wire net346;
wire net4;
wire net43;
wire net361;
wire net115;
wire net670;
wire in18;
wire net27;
wire net34;
wire net216;
wire net187;
wire in13;
wire net586;
wire net533;
wire net796;
wire net32;
wire net125;
wire net19;
wire in15;
wire net727;
wire net163;
wire in19;
wire net702;
wire net70;
wire net48;
wire net28;
wire net92;
wire net713;
wire net25;
wire out36;
wire net30;
wire in0;
wire net709;
wire net24;
wire out47;
wire net290;
wire net227;
wire net470;
wire in33;
wire net33;
wire net824;
wire net233;
wire net121;
wire net40;
wire in60;
wire net435;
wire net301;
wire net760;
wire net23;
wire net26;
wire net16;
wire net558;
wire in1;
wire net265;
wire in28;
wire net778;
wire net22;
wire net263;
wire net5;
wire net206;
wire in58;
wire in61;
wire net757;
wire in56;
wire net733;
wire net171;
wire in23;
wire out4;
wire net42;
wire net91;
wire in57;
wire net281;
wire net54;
wire net313;
wire in54;
wire in53;
wire net138;
wire net145;
wire net211;
wire in35;
wire in34;
wire net593;
wire in45;
wire net393;
wire net256;
wire net87;
wire net181;
wire net7;
wire net574;
wire net455;
wire net191;
wire out46;
wire in44;
wire in32;
wire net47;
wire net12;
wire in27;
wire in9;
wire net654;
wire net723;
wire net611;
wire net515;
wire net362;
wire in16;
wire net35;
wire net220;
wire in22;
wire net68;
wire in14;
wire net529;
wire in21;
wire net57;
wire net480;
wire net86;
wire net317;
wire in51;
wire net93;
wire in47;
wire in2;
wire net718;
wire net658;
wire net105;
wire in11;
wire net51;
wire in36;
wire net536;
wire net37;
wire net36;
wire net95;
wire net146;
wire net734;
wire net251;
wire net768;
wire net11;
wire net352;
wire net845;
wire net307;
wire net394;
wire net314;
wire in3;
sky130_fd_sc_hd__mux4_2 c62(
.A0(in50),
.A1(in57),
.A2(in61),
.A3(in59),
.S0(in58),
.S1(in25),
.X(net0)
);

sky130_fd_sc_hd__mux4_2 c63(
.A0(net0),
.A1(in49),
.A2(in45),
.A3(in44),
.S0(in56),
.S1(in50),
.X(net1)
);

sky130_fd_sc_hd__mux4_4 c64(
.A0(net3),
.A1(in54),
.A2(in53),
.A3(in50),
.S0(in47),
.S1(in45),
.X(net2)
);

sky130_fd_sc_hd__mux4_1 c65(
.A0(in13),
.A1(in29),
.A2(in25),
.A3(in26),
.S0(in35),
.S1(in36),
.X(net3)
);

sky130_fd_sc_hd__nand3_2 c66(
.A(in44),
.B(in59),
.C(in0),
.Y(net4)
);

sky130_fd_sc_hd__or4bb_4 c67(
.A(in47),
.B(in51),
.C_N(in31),
.D_N(in52),
.X(net5)
);

sky130_fd_sc_hd__nand3_4 c68(
.A(in52),
.B(net2),
.C(net5),
.Y(net6)
);

sky130_fd_sc_hd__o2111a_2 c69(
.A1(in56),
.A2(in0),
.B1(in61),
.C1(in45),
.D1(in48),
.X(net7)
);

sky130_fd_sc_hd__or3_4 c70(
.A(in34),
.B(net3),
.C(net7),
.X(net8)
);

sky130_fd_sc_hd__nand3_4 c71(
.A(net8),
.B(in59),
.C(in61),
.Y(net9)
);

sky130_fd_sc_hd__nand3_2 c72(
.A(in59),
.B(net9),
.C(net8),
.Y(net10)
);

sky130_fd_sc_hd__a2111oi_1 c73(
.A1(in60),
.A2(net10),
.B1(in61),
.C1(net5),
.D1(in0),
.Y(net11)
);

sky130_fd_sc_hd__o2111ai_1 c74(
.A1(net11),
.A2(in36),
.B1(net10),
.C1(in61),
.D1(net5),
.Y(net12)
);

sky130_fd_sc_hd__a2111oi_1 c75(
.A1(net9),
.A2(in60),
.B1(net11),
.C1(net10),
.D1(in25),
.Y(net13)
);

sky130_fd_sc_hd__a2111o_1 c76(
.A1(net5),
.A2(in52),
.B1(net13),
.C1(in44),
.D1(net2),
.X(net14)
);

sky130_fd_sc_hd__o2111ai_1 c77(
.A1(net9),
.A2(net11),
.B1(in25),
.C1(in20),
.D1(net8),
.Y(net15)
);

sky130_fd_sc_hd__mux4_2 c78(
.A0(net2),
.A1(net9),
.A2(in59),
.A3(net7),
.S0(net12),
.S1(net11),
.X(net16)
);

sky130_fd_sc_hd__or3b_1 c79(
.A(in49),
.B(net13),
.C_N(net10),
.X(net17)
);

sky130_fd_sc_hd__and3_2 c80(
.A(net12),
.B(net6),
.C(net10),
.X(net18)
);

sky130_fd_sc_hd__o2111a_4 c81(
.A1(in28),
.A2(net17),
.B1(net5),
.C1(net14),
.D1(in48),
.X(net19)
);

sky130_fd_sc_hd__nor3_1 c82(
.A(net16),
.B(net14),
.C(in54),
.Y(net20)
);

sky130_fd_sc_hd__and3_1 c83(
.A(net15),
.B(net8),
.C(net20),
.X(net21)
);

sky130_fd_sc_hd__a2111o_4 c84(
.A1(net21),
.A2(net16),
.B1(net14),
.C1(net17),
.D1(net8),
.X(net22)
);

sky130_fd_sc_hd__mux4_1 c85(
.A0(net22),
.A1(net21),
.A2(net10),
.A3(net17),
.S0(net5),
.S1(net20),
.X(net23)
);

sky130_fd_sc_hd__mux4_4 c86(
.A0(net18),
.A1(net22),
.A2(net23),
.A3(net21),
.S0(in37),
.S1(net19),
.X(net24)
);

sky130_fd_sc_hd__mux4_4 c87(
.A0(net24),
.A1(net18),
.A2(net17),
.A3(in29),
.S0(net23),
.S1(net22),
.X(net25)
);

sky130_fd_sc_hd__or3b_2 c88(
.A(net13),
.B(in7),
.C_N(in0),
.X(out29)
);

sky130_fd_sc_hd__or3_4 c89(
.A(in58),
.B(net5),
.C(in36),
.X(net26)
);

sky130_fd_sc_hd__or3_1 c90(
.A(net8),
.B(in45),
.C(in2),
.X(net27)
);

sky130_fd_sc_hd__nand3b_4 c91(
.A_N(net26),
.B(in31),
.C(net18),
.Y(net28)
);

sky130_fd_sc_hd__and3b_1 c92(
.A_N(net25),
.B(net22),
.C(net27),
.X(net29)
);

sky130_fd_sc_hd__nand3_4 c93(
.A(in7),
.B(net25),
.C(net28),
.Y(net30)
);

sky130_fd_sc_hd__or3_2 c94(
.A(net28),
.B(in37),
.C(net30),
.X(net31)
);

sky130_fd_sc_hd__or3b_2 c95(
.A(in20),
.B(net29),
.C_N(in51),
.X(net32)
);

sky130_fd_sc_hd__clkinv_1 c96(
.A(net665),
.Y(net33)
);

sky130_fd_sc_hd__buf_2 c97(
.A(net665),
.X(net34)
);

sky130_fd_sc_hd__sdfrbp_1 c98(
.D(net27),
.RESET_B(net31),
.SCD(net30),
.SCE(net34),
.CLK(clk),
.Q(net36),
.Q_N(net35)
);

sky130_fd_sc_hd__or4bb_2 c99(
.A(in54),
.B(in61),
.C_N(in48),
.D_N(net34),
.X(net37)
);

sky130_fd_sc_hd__a2111oi_1 c100(
.A1(net28),
.A2(net15),
.B1(net26),
.C1(net35),
.D1(net34),
.Y(net38)
);

sky130_fd_sc_hd__nor3_4 c101(
.A(net38),
.B(net29),
.C(net34),
.Y(net39)
);

sky130_fd_sc_hd__sdfbbn_1 c102(
.D(net37),
.RESET_B(net39),
.SCD(net38),
.SCE(net17),
.SET_B(net34),
.CLK_N(clk),
.Q(out55),
.Q_N(net40)
);

sky130_fd_sc_hd__a2111o_1 c103(
.A1(net39),
.A2(net31),
.B1(out55),
.C1(net38),
.D1(net34),
.X(net41)
);

sky130_fd_sc_hd__a2111oi_4 c104(
.A1(net33),
.A2(out55),
.B1(net38),
.C1(out29),
.D1(in20),
.Y(net42)
);

sky130_fd_sc_hd__mux4_1 c105(
.A0(net32),
.A1(net4),
.A2(net39),
.A3(net40),
.S0(net33),
.S1(in36),
.X(net43)
);

sky130_fd_sc_hd__sdfbbn_2 c106(
.D(net31),
.RESET_B(out55),
.SCD(net42),
.SCE(net38),
.SET_B(net37),
.CLK_N(clk),
.Q(net45),
.Q_N(net44)
);

sky130_fd_sc_hd__a2111oi_2 c107(
.A1(in45),
.A2(out55),
.B1(net34),
.C1(net702),
.D1(net755),
.Y(net46)
);

sky130_fd_sc_hd__mux4_4 c108(
.A0(net45),
.A1(out55),
.A2(net46),
.A3(net29),
.S0(net34),
.S1(net702),
.X(out53)
);

sky130_fd_sc_hd__mux4_1 c109(
.A0(net42),
.A1(net46),
.A2(out53),
.A3(net44),
.S0(net40),
.S1(net702),
.X(net47)
);

sky130_fd_sc_hd__buf_8 c110(
.A(net743),
.X(net48)
);

sky130_fd_sc_hd__dlygate4sd3_1 c111(
.A(net743),
.X(net49)
);

sky130_fd_sc_hd__nand3b_4 c112(
.A_N(net22),
.B(net48),
.C(net40),
.Y(net50)
);

sky130_fd_sc_hd__dfbbn_1 c113(
.D(net48),
.RESET_B(out53),
.SET_B(out29),
.CLK_N(clk),
.Q(out28),
.Q_N(net51)
);

sky130_fd_sc_hd__nand3_2 c114(
.A(net15),
.B(net48),
.C(in36),
.Y(out45)
);

sky130_fd_sc_hd__or3b_4 c115(
.A(in13),
.B(net48),
.C_N(net49),
.X(net52)
);

sky130_fd_sc_hd__nor3_2 c116(
.A(net45),
.B(net5),
.C(net52),
.Y(out46)
);

sky130_fd_sc_hd__mux4_1 c117(
.A0(net32),
.A1(in36),
.A2(out28),
.A3(out46),
.S0(net48),
.S1(net31),
.X(net53)
);

sky130_fd_sc_hd__or4bb_1 c118(
.A(net5),
.B(out46),
.C_N(net51),
.D_N(net756),
.X(net54)
);

sky130_fd_sc_hd__o2111a_4 c119(
.A1(out46),
.A2(in46),
.B1(net5),
.C1(net48),
.D1(out36),
.X(out51)
);

sky130_fd_sc_hd__o2111a_2 c120(
.A1(net50),
.A2(net48),
.B1(in13),
.C1(out46),
.D1(out28),
.X(net55)
);

sky130_fd_sc_hd__nor3_1 c121(
.A(net54),
.B(out46),
.C(out29),
.Y(net56)
);

sky130_fd_sc_hd__o2111ai_4 c122(
.A1(net52),
.A2(net5),
.B1(out28),
.C1(net56),
.D1(net48),
.Y(net57)
);

sky130_fd_sc_hd__or3b_1 c123(
.A(net48),
.B(out46),
.C_N(net17),
.X(net58)
);

sky130_fd_sc_hd__mux4_2 c124(
.A0(net55),
.A1(net32),
.A2(net52),
.A3(net56),
.S0(net54),
.S1(out46),
.X(net59)
);

sky130_fd_sc_hd__o2111ai_1 c125(
.A1(net10),
.A2(out28),
.B1(net48),
.C1(out46),
.D1(net50),
.Y(net60)
);

sky130_fd_sc_hd__or4bb_4 c126(
.A(net60),
.B(out46),
.C_N(in0),
.D_N(net17),
.X(net61)
);

sky130_fd_sc_hd__mux4_4 c127(
.A0(net57),
.A1(net22),
.A2(net15),
.A3(net48),
.S0(net60),
.S1(in46),
.X(net62)
);

sky130_fd_sc_hd__o2111a_1 c128(
.A1(net58),
.A2(net51),
.B1(net62),
.C1(net57),
.D1(out53),
.X(net63)
);

sky130_fd_sc_hd__sdfbbp_1 c129(
.D(net61),
.RESET_B(net62),
.SCD(net31),
.SCE(out46),
.SET_B(net744),
.CLK(clk),
.Q(net65),
.Q_N(net64)
);

sky130_fd_sc_hd__or4bb_1 c130(
.A(net56),
.B(net62),
.C_N(out46),
.D_N(net64),
.X(net66)
);

sky130_fd_sc_hd__mux4_2 c131(
.A0(net66),
.A1(in46),
.A2(net62),
.A3(out51),
.S0(net60),
.S1(out46),
.X(net67)
);

sky130_fd_sc_hd__or3_4 c132(
.A(in6),
.B(in1),
.C(in0),
.X(net68)
);

sky130_fd_sc_hd__or3b_1 c133(
.A(in6),
.B(in8),
.C_N(net68),
.X(net69)
);

sky130_fd_sc_hd__a2111oi_2 c134(
.A1(in19),
.A2(in9),
.B1(net68),
.C1(in4),
.D1(in8),
.Y(net70)
);

sky130_fd_sc_hd__or3_2 c135(
.A(in5),
.B(in10),
.C(in0),
.X(net71)
);

sky130_fd_sc_hd__o2111ai_4 c136(
.A1(in11),
.A2(net69),
.B1(net71),
.C1(in0),
.D1(net70),
.Y(net72)
);

sky130_fd_sc_hd__a2111o_1 c137(
.A1(in12),
.A2(in0),
.B1(in3),
.C1(net70),
.D1(net72),
.X(net73)
);

sky130_fd_sc_hd__nor3_1 c138(
.A(net68),
.B(net69),
.C(net72),
.Y(net74)
);

sky130_fd_sc_hd__a2111o_1 c139(
.A1(net74),
.A2(in14),
.B1(in1),
.C1(net68),
.D1(in0),
.X(net75)
);

sky130_fd_sc_hd__or4bb_1 c140(
.A(net73),
.B(net69),
.C_N(in14),
.D_N(in0),
.X(net76)
);

sky130_fd_sc_hd__mux4_2 c141(
.A0(in10),
.A1(net71),
.A2(in16),
.A3(net76),
.S0(net74),
.S1(net72),
.X(net77)
);

sky130_fd_sc_hd__a2111o_2 c142(
.A1(in4),
.A2(net74),
.B1(in1),
.C1(net73),
.D1(in0),
.X(net78)
);

sky130_fd_sc_hd__a2111oi_0 c143(
.A1(net71),
.A2(net74),
.B1(in8),
.C1(net69),
.D1(in0),
.Y(net79)
);

sky130_fd_sc_hd__a2111oi_0 c144(
.A1(in1),
.A2(net72),
.B1(net70),
.C1(net68),
.D1(net74),
.Y(net80)
);

sky130_fd_sc_hd__o2111ai_2 c145(
.A1(net75),
.A2(net73),
.B1(net80),
.C1(net79),
.D1(net78),
.Y(net81)
);

sky130_fd_sc_hd__a2111oi_4 c146(
.A1(net79),
.A2(in15),
.B1(net78),
.C1(net74),
.D1(net81),
.Y(net82)
);

sky130_fd_sc_hd__o2111ai_1 c147(
.A1(in15),
.A2(in21),
.B1(net70),
.C1(in13),
.D1(net80),
.Y(net83)
);

sky130_fd_sc_hd__o2111a_4 c148(
.A1(in8),
.A2(net82),
.B1(net80),
.C1(in14),
.D1(in5),
.X(net84)
);

sky130_fd_sc_hd__mux4_4 c149(
.A0(net69),
.A1(net76),
.A2(net79),
.A3(net78),
.S0(net68),
.S1(net74),
.X(net85)
);

sky130_fd_sc_hd__a2111o_2 c150(
.A1(in9),
.A2(in19),
.B1(net68),
.C1(net78),
.D1(net80),
.X(net86)
);

sky130_fd_sc_hd__o2111ai_2 c151(
.A1(net86),
.A2(in12),
.B1(in0),
.C1(net81),
.D1(net78),
.Y(net87)
);

sky130_fd_sc_hd__mux4_2 c152(
.A0(net83),
.A1(net87),
.A2(net80),
.A3(net86),
.S0(net72),
.S1(net69),
.X(net88)
);

sky130_fd_sc_hd__mux4_2 c153(
.A0(net88),
.A1(in8),
.A2(net87),
.A3(net78),
.S0(net69),
.S1(net86),
.X(net89)
);

sky130_fd_sc_hd__o2111ai_4 c154(
.A1(in30),
.A2(net84),
.B1(net85),
.C1(in0),
.D1(in31),
.Y(net90)
);

sky130_fd_sc_hd__or4bb_1 c155(
.A(in21),
.B(in35),
.C_N(net90),
.D_N(net72),
.X(net91)
);

sky130_fd_sc_hd__o2111ai_4 c156(
.A1(in17),
.A2(net87),
.B1(net80),
.C1(in36),
.D1(in22),
.Y(net92)
);

sky130_fd_sc_hd__or4bb_2 c157(
.A(in40),
.B(in41),
.C_N(in4),
.D_N(in29),
.X(net93)
);

sky130_fd_sc_hd__mux4_4 c158(
.A0(in39),
.A1(in22),
.A2(net90),
.A3(net72),
.S0(net93),
.S1(in27),
.X(net94)
);

sky130_fd_sc_hd__mux4_4 c159(
.A0(net91),
.A1(net94),
.A2(net90),
.A3(net93),
.S0(net76),
.S1(net68),
.X(net95)
);

sky130_fd_sc_hd__a2111o_4 c160(
.A1(in24),
.A2(in26),
.B1(net92),
.C1(net68),
.D1(in42),
.X(net96)
);

sky130_fd_sc_hd__or4bb_2 c161(
.A(in18),
.B(in23),
.C_N(in32),
.D_N(net69),
.X(net97)
);

sky130_fd_sc_hd__or4bb_2 c162(
.A(net97),
.B(in26),
.C_N(in0),
.D_N(in24),
.X(net98)
);

sky130_fd_sc_hd__a2111oi_4 c163(
.A1(in36),
.A2(in23),
.B1(net80),
.C1(in4),
.D1(net98),
.Y(net99)
);

sky130_fd_sc_hd__a2111oi_4 c164(
.A1(net94),
.A2(net93),
.B1(net85),
.C1(net70),
.D1(in25),
.Y(net100)
);

sky130_fd_sc_hd__nand3_1 c165(
.A(net100),
.B(in24),
.C(net95),
.Y(net101)
);

sky130_fd_sc_hd__mux4_4 c166(
.A0(in43),
.A1(net97),
.A2(net92),
.A3(in4),
.S0(net94),
.S1(net100),
.X(net102)
);

sky130_fd_sc_hd__mux4_2 c167(
.A0(net102),
.A1(net100),
.A2(net91),
.A3(in26),
.S0(net87),
.S1(net80),
.X(net103)
);

sky130_fd_sc_hd__a2111oi_1 c168(
.A1(in3),
.A2(net91),
.B1(net101),
.C1(in36),
.D1(net96),
.Y(net104)
);

sky130_fd_sc_hd__mux4_4 c169(
.A0(net101),
.A1(in18),
.A2(in26),
.A3(net98),
.S0(net104),
.S1(in39),
.X(net105)
);

sky130_fd_sc_hd__mux4_2 c170(
.A0(net87),
.A1(net102),
.A2(net103),
.A3(net94),
.S0(in39),
.S1(net101),
.X(net106)
);

sky130_fd_sc_hd__a2111oi_2 c171(
.A1(net92),
.A2(net106),
.B1(net104),
.C1(net99),
.D1(net101),
.Y(net107)
);

sky130_fd_sc_hd__mux4_2 c172(
.A0(in22),
.A1(net105),
.A2(net99),
.A3(net106),
.S0(net94),
.S1(net107),
.X(net108)
);

sky130_fd_sc_hd__mux4_4 c173(
.A0(net103),
.A1(net105),
.A2(net102),
.A3(net107),
.S0(net96),
.S1(net106),
.X(net109)
);

sky130_fd_sc_hd__mux4_2 c174(
.A0(net106),
.A1(net68),
.A2(net90),
.A3(net107),
.S0(net698),
.S1(net758),
.X(net110)
);

sky130_fd_sc_hd__mux4_1 c175(
.A0(net93),
.A1(net101),
.A2(net103),
.A3(net107),
.S0(net98),
.S1(net105),
.X(net111)
);

sky130_fd_sc_hd__or3_4 c176(
.A(net1),
.B(net99),
.C(in32),
.X(net112)
);

sky130_fd_sc_hd__or4bb_2 c177(
.A(net72),
.B(net90),
.C_N(in48),
.D_N(net757),
.X(net113)
);

sky130_fd_sc_hd__or4bb_1 c178(
.A(in26),
.B(net107),
.C_N(net113),
.D_N(in53),
.X(net114)
);

sky130_fd_sc_hd__a2111o_2 c179(
.A1(net98),
.A2(net1),
.B1(in46),
.C1(in48),
.D1(net750),
.X(net115)
);

sky130_fd_sc_hd__mux4_4 c180(
.A0(in16),
.A1(net92),
.A2(in48),
.A3(net99),
.S0(net115),
.S1(net750),
.X(net116)
);

sky130_fd_sc_hd__mux4_1 c181(
.A0(in55),
.A1(in25),
.A2(net89),
.A3(in61),
.S0(net115),
.S1(net750),
.X(net117)
);

sky130_fd_sc_hd__or4bb_2 c182(
.A(net105),
.B(net98),
.C_N(net85),
.D_N(in0),
.X(net118)
);

sky130_fd_sc_hd__mux4_1 c183(
.A0(in4),
.A1(net115),
.A2(in61),
.A3(net112),
.S0(net92),
.S1(net750),
.X(net119)
);

sky130_fd_sc_hd__mux4_2 c184(
.A0(net119),
.A1(net116),
.A2(net118),
.A3(net115),
.S0(net117),
.S1(net70),
.X(net120)
);

sky130_fd_sc_hd__mux4_1 c185(
.A0(net89),
.A1(net112),
.A2(net3),
.A3(net106),
.S0(in55),
.S1(net119),
.X(net121)
);

sky130_fd_sc_hd__o2111ai_2 c186(
.A1(in32),
.A2(in4),
.B1(net99),
.C1(net77),
.D1(out5),
.Y(net122)
);

sky130_fd_sc_hd__or3_1 c187(
.A(net113),
.B(net112),
.C(in37),
.X(net123)
);

sky130_fd_sc_hd__mux4_1 c188(
.A0(in50),
.A1(net97),
.A2(net123),
.A3(in26),
.S0(net122),
.S1(out5),
.X(net124)
);

sky130_fd_sc_hd__o2111ai_2 c189(
.A1(net107),
.A2(net121),
.B1(in4),
.C1(net116),
.D1(net123),
.Y(net125)
);

sky130_fd_sc_hd__or4bb_1 c190(
.A(net123),
.B(net124),
.C_N(in25),
.D_N(net118),
.X(net126)
);

sky130_fd_sc_hd__mux4_1 c191(
.A0(net123),
.A1(net124),
.A2(net113),
.A3(net122),
.S0(net643),
.S1(out5),
.X(net127)
);

sky130_fd_sc_hd__o2111a_2 c192(
.A1(net116),
.A2(net117),
.B1(net127),
.C1(net112),
.D1(net643),
.X(net128)
);

sky130_fd_sc_hd__mux4_2 c193(
.A0(net123),
.A1(net124),
.A2(net119),
.A3(net97),
.S0(net643),
.S1(net750),
.X(net129)
);

sky130_fd_sc_hd__mux4_2 c194(
.A0(net122),
.A1(in50),
.A2(in31),
.A3(net117),
.S0(net127),
.S1(net644),
.X(net130)
);

sky130_fd_sc_hd__mux4_2 c195(
.A0(net128),
.A1(net95),
.A2(net129),
.A3(net106),
.S0(net123),
.S1(net124),
.X(net131)
);

sky130_fd_sc_hd__mux4_4 c196(
.A0(net121),
.A1(net131),
.A2(net129),
.A3(net119),
.S0(net105),
.S1(net643),
.X(net132)
);

sky130_fd_sc_hd__mux4_1 c197(
.A0(net130),
.A1(net129),
.A2(net128),
.A3(net118),
.S0(net116),
.X(net709)
);

sky130_fd_sc_hd__a2111oi_0 c198(
.A1(net20),
.A2(net14),
.B1(net0),
.C1(net130),
.D1(net70),
.Y(net134)
);

sky130_fd_sc_hd__mux4_4 c199(
.A0(net6),
.A1(net70),
.A2(in35),
.A3(net122),
.S0(in48),
.S1(net85),
.X(net135)
);

sky130_fd_sc_hd__a2111oi_1 c200(
.A1(in53),
.A2(net23),
.B1(net90),
.C1(net68),
.D1(net708),
.Y(net136)
);

sky130_fd_sc_hd__sdfbbn_1 c201(
.D(net134),
.RESET_B(net20),
.SCD(in37),
.SCE(net130),
.SET_B(in25),
.CLK_N(clk),
.Q(net138),
.Q_N(net137)
);

sky130_fd_sc_hd__mux4_2 c202(
.A0(net121),
.A1(in37),
.A2(net112),
.A3(net21),
.S0(net119),
.S1(in0),
.X(net139)
);

sky130_fd_sc_hd__a2111oi_4 c203(
.A1(in61),
.A2(net127),
.B1(net17),
.C1(net7),
.D1(net130),
.Y(net140)
);

sky130_fd_sc_hd__o2111a_2 c204(
.A1(net138),
.A2(in57),
.B1(net14),
.C1(net698),
.D1(net708),
.X(net141)
);

sky130_fd_sc_hd__mux4_1 c205(
.A0(in53),
.A1(net138),
.A2(net140),
.A3(net90),
.S0(net70),
.S1(net708),
.X(net142)
);

sky130_fd_sc_hd__a2111o_1 c206(
.A1(net23),
.A2(net121),
.B1(net138),
.C1(net106),
.D1(net136),
.X(net143)
);

sky130_fd_sc_hd__mux4_1 c207(
.A0(net140),
.A1(net119),
.A2(net98),
.A3(net137),
.S0(net705),
.S1(out5),
.X(net144)
);

sky130_fd_sc_hd__mux4_2 c208(
.A0(net136),
.A1(in53),
.A2(net21),
.A3(net20),
.S0(net744),
.S1(net759),
.X(net145)
);

sky130_fd_sc_hd__sdfbbn_2 c209(
.D(net127),
.RESET_B(net135),
.SCD(in57),
.SCE(net137),
.SET_B(net140),
.CLK_N(clk),
.Q(net147),
.Q_N(net146)
);

sky130_fd_sc_hd__mux4_1 c210(
.A0(net140),
.A1(in37),
.A2(net6),
.A3(net146),
.S0(net90),
.S1(net759),
.X(net148)
);

sky130_fd_sc_hd__a2111oi_1 c211(
.A1(net138),
.A2(net146),
.B1(net106),
.C1(net141),
.D1(net759),
.Y(net149)
);

sky130_fd_sc_hd__mux4_4 c212(
.A0(net135),
.A1(net130),
.A2(net12),
.A3(net140),
.S0(net743),
.S1(net759),
.X(net150)
);

sky130_fd_sc_hd__mux4_2 c213(
.A0(net145),
.A1(net149),
.A2(net137),
.A3(net92),
.S0(net122),
.S1(net708),
.X(net151)
);

sky130_fd_sc_hd__a2111oi_0 c214(
.A1(in25),
.A2(net6),
.B1(net145),
.C1(net705),
.D1(net743),
.Y(out31)
);

sky130_fd_sc_hd__o2111ai_2 c215(
.A1(net20),
.A2(in48),
.B1(out31),
.C1(net149),
.D1(net743),
.Y(net152)
);

sky130_fd_sc_hd__a2111oi_1 c216(
.A1(net141),
.A2(out31),
.B1(net7),
.C1(net14),
.D1(net744),
.Y(net153)
);

sky130_fd_sc_hd__mux4_4 c217(
.A0(net153),
.A1(net146),
.A2(out31),
.A3(net744),
.S0(out5),
.S1(net759),
.X(net154)
);

sky130_fd_sc_hd__mux4_2 c218(
.A0(net80),
.A1(net153),
.A2(net92),
.A3(net680),
.S0(net743),
.S1(net759),
.X(net155)
);

sky130_fd_sc_hd__mux4_4 c219(
.A0(net14),
.A1(net3),
.A2(net140),
.A3(net137),
.S0(net680),
.S1(net759),
.X(net156)
);

sky130_fd_sc_hd__mux4_2 c220(
.A0(net112),
.A1(net17),
.A2(net140),
.A3(out31),
.S0(net70),
.S1(out48),
.X(net157)
);

sky130_fd_sc_hd__mux4_2 c221(
.A0(net90),
.A1(net4),
.A2(net147),
.A3(net140),
.S0(net112),
.S1(net761),
.X(net158)
);

sky130_fd_sc_hd__mux4_1 c222(
.A0(net70),
.A1(net36),
.A2(in57),
.A3(net106),
.S0(net34),
.S1(net666),
.X(out12)
);

sky130_fd_sc_hd__mux4_4 c223(
.A0(net153),
.A1(net35),
.A2(out48),
.A3(net755),
.S0(out52),
.S1(net761),
.X(net159)
);

sky130_fd_sc_hd__mux4_1 c224(
.A0(out55),
.A1(net68),
.A2(net153),
.A3(net666),
.S0(net681),
.S1(net764),
.X(net160)
);

sky130_fd_sc_hd__mux4_2 c225(
.A0(net147),
.A1(out12),
.A2(net705),
.A3(out52),
.S0(net762),
.S1(net765),
.X(net161)
);

sky130_fd_sc_hd__mux4_2 c226(
.A0(out12),
.A1(net30),
.A2(net17),
.A3(net81),
.S0(net756),
.S1(net761),
.X(net162)
);

sky130_fd_sc_hd__mux4_4 c227(
.A0(net92),
.A1(in48),
.A2(out12),
.A3(net681),
.S0(net762),
.S1(net765),
.X(net163)
);

sky130_fd_sc_hd__mux4_1 c228(
.A0(net106),
.A1(net92),
.A2(net153),
.A3(net70),
.S0(net760),
.S1(net766),
.X(net164)
);

sky130_fd_sc_hd__mux4_1 c229(
.A0(net140),
.A1(in52),
.A2(out12),
.A3(net762),
.S0(net765),
.S1(net766),
.X(net165)
);

sky130_fd_sc_hd__mux4_2 c230(
.A0(net68),
.A1(net34),
.A2(net153),
.A3(net761),
.S0(net767),
.S1(net768),
.X(net166)
);

sky130_fd_sc_hd__mux4_4 c231(
.A0(in37),
.A1(in0),
.A2(net153),
.A3(net34),
.S0(net763),
.S1(net770),
.X(net167)
);

sky130_fd_sc_hd__mux4_4 c232(
.A0(in57),
.A1(net90),
.A2(net85),
.A3(net112),
.S0(net764),
.S1(net767),
.X(net168)
);

sky130_fd_sc_hd__mux4_4 c233(
.A0(net147),
.A1(net744),
.A2(net762),
.A3(out15),
.S0(net768),
.S1(net769),
.X(out58)
);

sky130_fd_sc_hd__mux4_1 c234(
.A0(net147),
.A1(net90),
.A2(in48),
.A3(out52),
.S0(net763),
.S1(net770),
.X(net169)
);

sky130_fd_sc_hd__mux4_1 c235(
.A0(net4),
.A1(net140),
.A2(out48),
.A3(net767),
.S0(net769),
.S1(net770),
.X(net170)
);

sky130_fd_sc_hd__mux4_2 c236(
.A0(net40),
.A1(in13),
.A2(net761),
.A3(net764),
.S0(net769),
.S1(net770),
.X(net171)
);

sky130_fd_sc_hd__mux4_1 c237(
.A0(net30),
.A1(net38),
.A2(net168),
.A3(net763),
.S0(net766),
.S1(net771),
.X(net172)
);

sky130_fd_sc_hd__mux4_2 c238(
.A0(net85),
.A1(net171),
.A2(net172),
.A3(net169),
.S0(out48),
.S1(net771),
.X(net173)
);

sky130_fd_sc_hd__mux4_4 c239(
.A0(net169),
.A1(net765),
.A2(net767),
.A3(net769),
.S0(net771),
.S1(net772),
.X(net174)
);

sky130_fd_sc_hd__mux4_1 c240(
.A0(net168),
.A1(net174),
.A2(net17),
.A3(out47),
.S0(out15),
.S1(net772),
.X(net175)
);

sky130_fd_sc_hd__mux4_4 c241(
.A0(net171),
.A1(net85),
.A2(net169),
.A3(net175),
.S0(net766),
.S1(net769),
.X(out44)
);

sky130_fd_sc_hd__mux4_2 c242(
.A0(net67),
.A1(net65),
.A2(net62),
.A3(net97),
.S0(in0),
.S1(net765),
.X(net176)
);

sky130_fd_sc_hd__mux4_2 c243(
.A0(net69),
.A1(in36),
.A2(out46),
.A3(in46),
.S0(out29),
.S1(out5),
.X(net177)
);

sky130_fd_sc_hd__mux4_4 c244(
.A0(net177),
.A1(out12),
.A2(net62),
.A3(out55),
.S0(net744),
.S1(net755),
.X(net178)
);

sky130_fd_sc_hd__mux4_1 c245(
.A0(net177),
.A1(net97),
.A2(net51),
.A3(net744),
.S0(out5),
.S1(out52),
.X(net179)
);

sky130_fd_sc_hd__mux4_2 c246(
.A0(net179),
.A1(net46),
.A2(out46),
.A3(in31),
.S0(net177),
.S1(out52),
.X(out22)
);

sky130_fd_sc_hd__mux4_4 c247(
.A0(net65),
.A1(net177),
.A2(out53),
.A3(out47),
.S0(out52),
.S1(net761),
.X(net180)
);

sky130_fd_sc_hd__mux4_2 c248(
.A0(net36),
.A1(net177),
.A2(net179),
.A3(net732),
.S0(net749),
.S1(net761),
.X(net181)
);

sky130_fd_sc_hd__mux4_4 c249(
.A0(net46),
.A1(net62),
.A2(in46),
.A3(net732),
.S0(net749),
.S1(out15),
.X(net182)
);

sky130_fd_sc_hd__mux4_1 c250(
.A0(net181),
.A1(net177),
.A2(net182),
.A3(net51),
.S0(out12),
.S1(out46),
.X(net183)
);

sky130_fd_sc_hd__mux4_1 c251(
.A0(net49),
.A1(in46),
.A2(net182),
.A3(net177),
.S0(net181),
.S1(out5),
.X(out57)
);

sky130_fd_sc_hd__mux4_4 c252(
.A0(net175),
.A1(in31),
.A2(net177),
.A3(out46),
.S0(net182),
.S1(net732),
.X(net184)
);

sky130_fd_sc_hd__mux4_1 c253(
.A0(in36),
.A1(net69),
.A2(net182),
.A3(net177),
.S0(net65),
.S1(net749),
.X(net185)
);

sky130_fd_sc_hd__mux4_1 c254(
.A0(net62),
.A1(net182),
.A2(net51),
.A3(net177),
.S0(net185),
.S1(out43),
.X(net186)
);

sky130_fd_sc_hd__mux4_4 c255(
.A0(net67),
.A1(net35),
.A2(net184),
.A3(out36),
.S0(net761),
.S1(net773),
.X(net187)
);

sky130_fd_sc_hd__mux4_2 c256(
.A0(net182),
.A1(in31),
.A2(net749),
.A3(out15),
.S0(out43),
.S1(net775),
.X(net188)
);

sky130_fd_sc_hd__mux4_4 c257(
.A0(net188),
.A1(net182),
.A2(net64),
.A3(net756),
.S0(net773),
.S1(net775),
.X(net189)
);

sky130_fd_sc_hd__mux4_1 c258(
.A0(net184),
.A1(net62),
.A2(net744),
.A3(out52),
.S0(out43),
.S1(net775),
.X(net190)
);

sky130_fd_sc_hd__mux4_4 c259(
.A0(out36),
.A1(net761),
.A2(net765),
.A3(out43),
.S0(net775),
.S1(net776),
.X(net191)
);

sky130_fd_sc_hd__mux4_1 c260(
.A0(net191),
.A1(net182),
.A2(net51),
.A3(net773),
.S0(net774),
.S1(net776),
.X(net192)
);

sky130_fd_sc_hd__mux4_1 c261(
.A0(net192),
.A1(net191),
.A2(out36),
.A3(net773),
.S0(net774),
.S1(net776),
.X(net193)
);

sky130_fd_sc_hd__mux4_4 c262(
.A0(net182),
.A1(net62),
.A2(out36),
.A3(net743),
.S0(net774),
.S1(net776),
.X(net194)
);

sky130_fd_sc_hd__mux4_4 c263(
.A0(net185),
.A1(net194),
.A2(net62),
.A3(net743),
.S0(net774),
.S1(net776),
.X(net195)
);

sky130_fd_sc_hd__and2_1 c264(
.A(net77),
.B(net72),
.X(net196)
);

sky130_fd_sc_hd__a2111o_1 c265(
.A1(net86),
.A2(in14),
.B1(net70),
.C1(in0),
.D1(net196),
.X(net197)
);

sky130_fd_sc_hd__nor2_4 c266(
.A(net70),
.B(net197),
.Y(net198)
);

sky130_fd_sc_hd__nand3_4 c267(
.A(net89),
.B(net198),
.C(net81),
.Y(net199)
);

sky130_fd_sc_hd__or3b_1 c268(
.A(net197),
.B(net83),
.C_N(net70),
.X(net200)
);

sky130_fd_sc_hd__and3b_2 c269(
.A_N(net199),
.B(in14),
.C(net200),
.X(net201)
);

sky130_fd_sc_hd__or4bb_1 c270(
.A(net199),
.B(net200),
.C_N(net196),
.D_N(net83),
.X(net202)
);

sky130_fd_sc_hd__and3_1 c271(
.A(net200),
.B(net202),
.C(net198),
.X(net203)
);

sky130_fd_sc_hd__nor3_4 c272(
.A(net198),
.B(net201),
.C(net202),
.Y(net204)
);

sky130_fd_sc_hd__and2_1 c273(
.A(net203),
.B(net204),
.X(net205)
);

sky130_fd_sc_hd__nand3b_1 c274(
.A_N(net205),
.B(net196),
.C(net204),
.Y(net206)
);

sky130_fd_sc_hd__and3b_1 c275(
.A_N(net205),
.B(net199),
.C(net204),
.X(net207)
);

sky130_fd_sc_hd__mux4_4 c276(
.A0(net71),
.A1(net206),
.A2(net205),
.A3(net196),
.S0(net70),
.S1(net72),
.X(net208)
);

sky130_fd_sc_hd__mux4_1 c277(
.A0(net79),
.A1(net207),
.A2(net201),
.A3(net205),
.S0(net199),
.S1(in2),
.X(net209)
);

sky130_fd_sc_hd__mux4_4 c278(
.A0(net208),
.A1(net196),
.A2(net202),
.A3(net204),
.S0(net209),
.S1(net70),
.X(net210)
);

sky130_fd_sc_hd__or4bb_2 c279(
.A(net201),
.B(net199),
.C_N(net207),
.D_N(net668),
.X(net211)
);

sky130_fd_sc_hd__sdfrbp_2 c280(
.D(net211),
.RESET_B(net205),
.SCD(net203),
.SCE(net668),
.CLK(clk),
.Q(net213),
.Q_N(net212)
);

sky130_fd_sc_hd__sdfbbp_1 c281(
.D(net207),
.RESET_B(net200),
.SCD(net211),
.SCE(in14),
.SET_B(net204),
.CLK(clk),
.Q(net215),
.Q_N(net214)
);

sky130_fd_sc_hd__o2111ai_2 c282(
.A1(net198),
.A2(net206),
.B1(net212),
.C1(net208),
.D1(net668),
.Y(net216)
);

sky130_fd_sc_hd__mux4_1 c283(
.A0(net213),
.A1(net75),
.A2(net206),
.A3(net198),
.S0(net196),
.S1(net674),
.X(net217)
);

sky130_fd_sc_hd__a2111o_1 c284(
.A1(net217),
.A2(net204),
.B1(net75),
.C1(net214),
.D1(net674),
.X(net218)
);

sky130_fd_sc_hd__mux4_4 c285(
.A0(net204),
.A1(net206),
.A2(net217),
.A3(net208),
.S0(net668),
.S1(net674),
.X(net219)
);

sky130_fd_sc_hd__or4bb_1 c286(
.A(in23),
.B(net78),
.C_N(in35),
.D_N(net777),
.X(net220)
);

sky130_fd_sc_hd__and3_4 c287(
.A(net78),
.B(net81),
.C(net95),
.X(net221)
);

sky130_fd_sc_hd__nand3b_4 c288(
.A_N(net96),
.B(net72),
.C(net698),
.Y(net222)
);

sky130_fd_sc_hd__or4bb_4 c289(
.A(net206),
.B(net95),
.C_N(net196),
.D_N(in0),
.X(net223)
);

sky130_fd_sc_hd__or4bb_1 c290(
.A(net220),
.B(net78),
.C_N(in27),
.D_N(net81),
.X(net224)
);

sky130_fd_sc_hd__or3b_2 c291(
.A(net96),
.B(net84),
.C_N(net222),
.X(net225)
);

sky130_fd_sc_hd__mux4_1 c292(
.A0(net225),
.A1(net223),
.A2(net222),
.A3(net209),
.S0(net78),
.S1(net96),
.X(net226)
);

sky130_fd_sc_hd__mux4_2 c293(
.A0(net224),
.A1(net222),
.A2(net223),
.A3(in23),
.S0(net698),
.S1(net777),
.X(net227)
);

sky130_fd_sc_hd__and3b_4 c294(
.A_N(net225),
.B(net674),
.C(out1),
.X(net228)
);

sky130_fd_sc_hd__nand3b_4 c295(
.A_N(net657),
.B(net668),
.C(out1),
.Y(net229)
);

sky130_fd_sc_hd__or4bb_2 c296(
.A(in38),
.B(net221),
.C_N(net202),
.D_N(net98),
.X(net230)
);

sky130_fd_sc_hd__nand3b_1 c297(
.A_N(net224),
.B(net230),
.C(net668),
.Y(net231)
);

sky130_fd_sc_hd__mux4_4 c298(
.A0(net230),
.A1(net224),
.A2(in35),
.A3(net203),
.S0(in27),
.S1(out1),
.X(net232)
);

sky130_fd_sc_hd__mux4_4 c299(
.A0(net223),
.A1(net98),
.A2(net232),
.A3(net222),
.X(net233),
.S1(net757)
);

sky130_fd_sc_hd__nand3b_2 c300(
.A_N(net72),
.B(net228),
.C(net668),
.Y(net234)
);

sky130_fd_sc_hd__or3b_1 c301(
.A(net232),
.B(net657),
.C_N(net698),
.X(out61)
);

sky130_fd_sc_hd__mux4_2 c302(
.A0(in33),
.A1(net232),
.A2(out61),
.A3(in4),
.S0(net96),
.S1(net657),
.X(net235)
);

sky130_fd_sc_hd__mux4_2 c303(
.A0(net89),
.A1(net223),
.A2(net97),
.A3(in31),
.S0(in0),
.S1(net778),
.X(net236)
);

sky130_fd_sc_hd__mux4_4 c304(
.A0(net221),
.A1(net96),
.A2(net657),
.A3(net668),
.S0(net674),
.S1(net698),
.X(net237)
);

sky130_fd_sc_hd__mux4_2 c305(
.A0(net234),
.A1(net96),
.A2(net228),
.A3(net673),
.S0(net698),
.S1(net778),
.X(net238)
);

sky130_fd_sc_hd__mux4_1 c306(
.A0(net234),
.A1(in41),
.A2(net96),
.A3(net223),
.S0(net232),
.S1(net673),
.X(net239)
);

sky130_fd_sc_hd__mux4_2 c307(
.A0(net229),
.A1(net224),
.A2(net202),
.A3(net232),
.S0(net230),
.S1(net673),
.X(net240)
);

sky130_fd_sc_hd__clkinv_8 c308(
.A(net738),
.Y(out38)
);

sky130_fd_sc_hd__nor3_2 c309(
.A(net117),
.B(net221),
.C(out5),
.Y(net241)
);

sky130_fd_sc_hd__a2111oi_4 c310(
.A1(net241),
.A2(in42),
.B1(net644),
.C1(net657),
.D1(net709),
.Y(net242)
);

sky130_fd_sc_hd__buf_12 c311(
.A(net738),
.X(net243)
);

sky130_fd_sc_hd__mux4_1 c312(
.A0(net84),
.A1(net241),
.A2(out38),
.A3(net72),
.S0(out61),
.S1(net709),
.X(net244)
);

sky130_fd_sc_hd__a2111oi_2 c313(
.A1(net221),
.A2(in52),
.B1(net76),
.C1(net644),
.D1(net780),
.Y(net245)
);

sky130_fd_sc_hd__a2111o_1 c314(
.A1(net129),
.A2(net245),
.B1(net99),
.C1(net778),
.D1(net780),
.X(net246)
);

sky130_fd_sc_hd__buf_2 c315(
.A(net672),
.X(net247)
);

sky130_fd_sc_hd__mux4_2 c316(
.A0(in42),
.A1(net245),
.A2(net117),
.A3(net246),
.S0(net131),
.S1(net95),
.X(net248)
);

sky130_fd_sc_hd__clkinv_4 c317(
.A(net672),
.Y(net249)
);

sky130_fd_sc_hd__mux4_2 c318(
.A0(net95),
.A1(out38),
.A2(net673),
.A3(net757),
.S0(net779),
.S1(net782),
.X(net250)
);

sky130_fd_sc_hd__mux4_2 c319(
.A0(net241),
.A1(net0),
.A2(net129),
.A3(in61),
.S0(net758),
.S1(net780),
.X(net251)
);

sky130_fd_sc_hd__mux4_2 c320(
.A0(net240),
.A1(net124),
.A2(net251),
.A3(in48),
.S0(net245),
.S1(net777),
.X(net252)
);

sky130_fd_sc_hd__mux4_2 c321(
.A0(in35),
.A1(net247),
.A2(net250),
.A3(net251),
.S0(net673),
.S1(net709),
.X(net253)
);

sky130_fd_sc_hd__sdfbbn_1 c322(
.D(net253),
.RESET_B(net246),
.SCD(net249),
.SCE(in0),
.SET_B(net750),
.CLK_N(clk),
.Q(net255),
.Q_N(net254)
);

sky130_fd_sc_hd__mux4_1 c323(
.A0(net118),
.A1(net255),
.A2(net241),
.A3(net251),
.S0(in31),
.S1(net215),
.X(net256)
);

sky130_fd_sc_hd__mux4_4 c324(
.A0(net99),
.A1(net255),
.A2(net251),
.A3(net242),
.S0(in48),
.S1(net698),
.X(net257)
);

sky130_fd_sc_hd__o2111ai_2 c325(
.A1(net240),
.A2(net255),
.B1(net209),
.C1(net750),
.D1(net777),
.Y(net258)
);

sky130_fd_sc_hd__mux4_2 c326(
.A0(net253),
.A1(net254),
.A2(net0),
.A3(net734),
.S0(net780),
.S1(net782),
.X(net259)
);

sky130_fd_sc_hd__mux4_1 c327(
.A0(net131),
.A1(net255),
.A2(net129),
.A3(net251),
.S0(net257),
.S1(out7),
.X(net260)
);

sky130_fd_sc_hd__a2111oi_2 c328(
.A1(net246),
.A2(in29),
.B1(net128),
.C1(net254),
.D1(net750),
.Y(net261)
);

sky130_fd_sc_hd__mux4_1 c329(
.A0(net261),
.A1(net128),
.A2(net254),
.A3(net657),
.S0(net750),
.S1(net783),
.X(net262)
);

sky130_fd_sc_hd__mux4_1 c330(
.A0(net221),
.A1(net7),
.A2(net153),
.A3(net98),
.S0(net760),
.S1(net777),
.X(net263)
);

sky130_fd_sc_hd__mux4_1 c331(
.A0(net251),
.A1(net249),
.A2(net149),
.A3(net760),
.S0(net779),
.S1(net782),
.X(net264)
);

sky130_fd_sc_hd__mux4_1 c332(
.A0(net21),
.A1(net251),
.A2(net149),
.A3(net138),
.S0(net209),
.S1(net786),
.X(net265)
);

sky130_fd_sc_hd__mux4_1 c333(
.A0(net149),
.A1(net119),
.A2(net221),
.A3(net124),
.X(net266),
.S1(net781)
);

sky130_fd_sc_hd__mux4_1 c334(
.A0(in41),
.A1(net70),
.A2(net137),
.A3(net153),
.S0(out52),
.S1(net780),
.X(net267)
);

sky130_fd_sc_hd__mux4_4 c335(
.A0(net128),
.A1(net130),
.A2(net153),
.A3(net237),
.S0(out52),
.S1(net788),
.X(net268)
);

sky130_fd_sc_hd__mux4_1 c336(
.A0(net0),
.A1(net149),
.A2(net21),
.A3(in0),
.S0(net781),
.S1(net788),
.X(net269)
);

sky130_fd_sc_hd__mux4_4 c337(
.A0(net12),
.A1(net18),
.A2(in46),
.A3(net149),
.S0(net746),
.S1(net777),
.X(net270)
);

sky130_fd_sc_hd__mux4_2 c338(
.A0(net3),
.A1(out61),
.A2(net204),
.A3(net746),
.S0(net786),
.S1(net790),
.X(net271)
);

sky130_fd_sc_hd__a2111o_1 c339(
.A1(net130),
.A2(net221),
.B1(net740),
.C1(net788),
.D1(net789),
.X(net272)
);

sky130_fd_sc_hd__mux4_4 c340(
.A0(net250),
.A1(net760),
.A2(net780),
.A3(net784),
.S0(net788),
.S1(net790),
.X(net273)
);

sky130_fd_sc_hd__mux4_1 c341(
.A0(net272),
.A1(net250),
.A2(net21),
.A3(net661),
.S0(net746),
.S1(net779),
.X(net274)
);

sky130_fd_sc_hd__mux4_2 c342(
.A0(net273),
.A1(net130),
.A2(net247),
.A3(net661),
.S0(net781),
.S1(net785),
.X(net275)
);

sky130_fd_sc_hd__mux4_1 c343(
.A0(net7),
.A1(net149),
.A2(net662),
.A3(net777),
.S0(net786),
.S1(net790),
.X(net276)
);

sky130_fd_sc_hd__mux4_2 c344(
.A0(net273),
.A1(out61),
.A2(net115),
.A3(net275),
.S0(net746),
.S1(out56),
.X(net277)
);

sky130_fd_sc_hd__mux4_2 c345(
.A0(net273),
.A1(net153),
.A2(in29),
.A3(in0),
.S0(net788),
.S1(net794),
.X(net278)
);

sky130_fd_sc_hd__mux4_1 c346(
.A0(net272),
.A1(net119),
.A2(net733),
.A3(net739),
.S0(net780),
.S1(net794),
.X(net279)
);

sky130_fd_sc_hd__mux4_2 c347(
.A0(net245),
.A1(net272),
.A2(net7),
.A3(net249),
.S0(net750),
.S1(out56),
.X(net280)
);

sky130_fd_sc_hd__mux4_1 c348(
.A0(net727),
.A1(net733),
.A2(net790),
.A3(net791),
.S0(net794),
.S1(net795),
.X(net281)
);

sky130_fd_sc_hd__mux4_1 c349(
.A0(out31),
.A1(net733),
.A2(net739),
.A3(net786),
.S0(net788),
.S1(net795),
.X(net282)
);

sky130_fd_sc_hd__mux4_4 c350(
.A0(net282),
.A1(net12),
.A2(net281),
.A3(net727),
.S0(net787),
.S1(net794),
.X(net283)
);

sky130_fd_sc_hd__mux4_4 c351(
.A0(net281),
.A1(net4),
.A2(net662),
.A3(net727),
.S0(net733),
.S1(net795),
.X(net284)
);

sky130_fd_sc_hd__mux4_4 c352(
.A0(net4),
.A1(net70),
.A2(net119),
.A3(net40),
.S0(in13),
.S1(net115),
.X(net285)
);

sky130_fd_sc_hd__mux4_1 c353(
.A0(net275),
.A1(net70),
.A2(net740),
.A3(net760),
.S0(net765),
.S1(net769),
.X(net286)
);

sky130_fd_sc_hd__mux4_1 c354(
.A0(net98),
.A1(net282),
.A2(net760),
.A3(net782),
.S0(net788),
.S1(net791),
.X(net287)
);

sky130_fd_sc_hd__sdfbbn_2 c355(
.D(out53),
.RESET_B(net740),
.SCD(net765),
.SCE(net772),
.SET_B(net786),
.CLK_N(clk),
.Q(net289),
.Q_N(net288)
);

sky130_fd_sc_hd__mux4_1 c356(
.A0(net40),
.A1(in52),
.A2(out5),
.A3(net771),
.S0(net782),
.S1(net786),
.X(out16)
);

sky130_fd_sc_hd__mux4_2 c357(
.A0(net282),
.A1(net209),
.A2(net249),
.A3(net34),
.S0(net772),
.S1(net796),
.X(net290)
);

sky130_fd_sc_hd__mux4_4 c358(
.A0(net285),
.A1(net77),
.A2(net282),
.A3(net765),
.S0(net770),
.S1(net791),
.X(net291)
);

sky130_fd_sc_hd__mux4_4 c359(
.A0(net289),
.A1(out16),
.A2(net725),
.A3(net740),
.S0(net768),
.S1(net786),
.X(out25)
);

sky130_fd_sc_hd__mux4_2 c360(
.A0(net247),
.A1(net213),
.A2(net70),
.A3(net288),
.S0(net745),
.S1(net765),
.X(net292)
);

sky130_fd_sc_hd__o2111ai_2 c361(
.A1(net292),
.A2(net275),
.B1(in2),
.C1(net40),
.D1(net17),
.Y(net293)
);

sky130_fd_sc_hd__o2111ai_2 c362(
.A1(net289),
.A2(net292),
.B1(out25),
.C1(net284),
.D1(net282),
.Y(net294)
);

sky130_fd_sc_hd__sdfbbp_1 c363(
.D(net153),
.RESET_B(out44),
.SCD(out61),
.SCE(out49),
.SET_B(net779),
.CLK(clk),
.Q(net296),
.Q_N(net295)
);

sky130_fd_sc_hd__mux4_1 c364(
.A0(net292),
.A1(net705),
.A2(out48),
.A3(net745),
.S0(net772),
.S1(net787),
.X(net297)
);

sky130_fd_sc_hd__mux4_1 c365(
.A0(net34),
.A1(out16),
.A2(net153),
.A3(net668),
.S0(net745),
.S1(net762),
.X(net298)
);

sky130_fd_sc_hd__mux4_2 c366(
.A0(net172),
.A1(in48),
.A2(net34),
.A3(out31),
.S0(net288),
.S1(out48),
.X(net299)
);

sky130_fd_sc_hd__mux4_2 c367(
.A0(net174),
.A1(net296),
.A2(net284),
.A3(net34),
.S0(net734),
.S1(net797),
.X(net300)
);

sky130_fd_sc_hd__mux4_4 c368(
.A0(net122),
.A1(in46),
.A2(net4),
.A3(net212),
.S0(net300),
.S1(net797),
.X(out32)
);

sky130_fd_sc_hd__mux4_2 c369(
.A0(in2),
.A1(net153),
.A2(net300),
.A3(net292),
.S0(net745),
.S1(net796),
.X(net301)
);

sky130_fd_sc_hd__mux4_4 c370(
.A0(net297),
.A1(net292),
.A2(net34),
.A3(out48),
.S0(net772),
.S1(net797),
.X(net302)
);

sky130_fd_sc_hd__mux4_1 c371(
.A0(net296),
.A1(net302),
.A2(net734),
.A3(net768),
.S0(net781),
.S1(net798),
.X(net303)
);

sky130_fd_sc_hd__mux4_4 c372(
.A0(net275),
.A1(net115),
.A2(net303),
.A3(in61),
.S0(out31),
.S1(net797),
.X(net304)
);

sky130_fd_sc_hd__mux4_2 c373(
.A0(net295),
.A1(out32),
.A2(net705),
.A3(net725),
.S0(net796),
.S1(net797),
.X(out50)
);

sky130_fd_sc_hd__mux4_1 c392(
.A0(out28),
.A1(out58),
.A2(out51),
.A3(out57),
.S0(out47),
.S1(net779),
.X(net305)
);

sky130_fd_sc_hd__mux4_4 c393(
.A0(net36),
.A1(net215),
.A2(out46),
.A3(out54),
.S0(net702),
.S1(out5),
.X(out60)
);

sky130_fd_sc_hd__mux4_1 c394(
.A0(net188),
.A1(out60),
.A2(out22),
.X(net306),
.S0(net702),
.S1(net779)
);

sky130_fd_sc_hd__o2111a_1 c395(
.A1(net17),
.A2(out60),
.B1(out54),
.C1(net702),
.D1(net779),
.X(out27)
);

sky130_fd_sc_hd__or2b_1 c396(
.A(net197),
.B_N(in13),
.X(net307)
);

sky130_fd_sc_hd__inv_6 c397(
.A(net675),
.Y(net308)
);

sky130_fd_sc_hd__clkbuf_2 c398(
.A(net675),
.X(net309)
);

sky130_fd_sc_hd__or3b_1 c399(
.A(net309),
.B(net197),
.C_N(net72),
.X(net310)
);

sky130_fd_sc_hd__and2b_2 c400(
.A_N(net310),
.B(net196),
.X(net311)
);

sky130_fd_sc_hd__and3b_2 c401(
.A_N(net73),
.B(in14),
.C(net311),
.X(net312)
);

sky130_fd_sc_hd__a2111oi_4 c402(
.A1(net312),
.A2(net77),
.B1(net211),
.C1(net72),
.D1(net203),
.Y(net313)
);

sky130_fd_sc_hd__mux4_4 c403(
.A0(net75),
.A1(net88),
.A2(net78),
.A3(net77),
.S0(net309),
.S1(in14),
.X(net314)
);

sky130_fd_sc_hd__or4bb_2 c404(
.A(net307),
.B(net312),
.C_N(net314),
.D_N(net202),
.X(net315)
);

sky130_fd_sc_hd__and3b_1 c405(
.A_N(net314),
.B(net307),
.C(net214),
.X(net316)
);

sky130_fd_sc_hd__or3_2 c406(
.A(net82),
.B(net311),
.C(net312),
.X(net317)
);

sky130_fd_sc_hd__nand3b_4 c407(
.A_N(net317),
.B(net308),
.C(in0),
.Y(net318)
);

sky130_fd_sc_hd__or4bb_4 c408(
.A(net314),
.B(net211),
.C_N(net317),
.D_N(net318),
.X(net319)
);

sky130_fd_sc_hd__nor3_1 c409(
.A(net318),
.B(net315),
.C(net649),
.Y(net320)
);

sky130_fd_sc_hd__o2111ai_4 c410(
.A1(net316),
.A2(net318),
.B1(net81),
.C1(net317),
.D1(net714),
.Y(net321)
);

sky130_fd_sc_hd__o2111a_2 c411(
.A1(net311),
.A2(net215),
.B1(net321),
.C1(net320),
.D1(in14),
.X(net322)
);

sky130_fd_sc_hd__mux4_4 c412(
.A0(net204),
.A1(net322),
.A2(net318),
.A3(net315),
.S0(net312),
.S1(net320),
.X(net323)
);

sky130_fd_sc_hd__o2111ai_2 c413(
.A1(net315),
.A2(net321),
.B1(net310),
.C1(net312),
.D1(net648),
.Y(net324)
);

sky130_fd_sc_hd__mux4_4 c414(
.A0(in14),
.A1(net324),
.A2(net318),
.A3(net310),
.S0(net312),
.S1(net649),
.X(net325)
);

sky130_fd_sc_hd__mux4_4 c415(
.A0(net322),
.A1(net197),
.A2(net312),
.A3(net320),
.S0(net316),
.S1(net714),
.X(net326)
);

sky130_fd_sc_hd__mux4_1 c416(
.A0(net317),
.A1(net324),
.A2(net318),
.A3(net204),
.S0(net320),
.S1(net648),
.X(net327)
);

sky130_fd_sc_hd__mux4_4 c417(
.A0(net312),
.A1(net72),
.A2(net318),
.A3(net714),
.S0(net800),
.S1(net803),
.X(net328)
);

sky130_fd_sc_hd__nor3_1 c418(
.A(net315),
.B(net200),
.C(net803),
.Y(net329)
);

sky130_fd_sc_hd__or3b_1 c419(
.A(net232),
.B(net778),
.C_N(net799),
.X(net330)
);

sky130_fd_sc_hd__nor3_4 c420(
.A(net238),
.B(net317),
.C(net232),
.Y(net331)
);

sky130_fd_sc_hd__nand3b_1 c421(
.A_N(net238),
.B(in13),
.C(net657),
.Y(net332)
);

sky130_fd_sc_hd__sdfrtn_1 c422(
.D(net308),
.RESET_B(net331),
.SCD(net657),
.SCE(net801),
.CLK_N(clk),
.Q(net333)
);

sky130_fd_sc_hd__sdfbbn_1 c423(
.D(net200),
.RESET_B(net332),
.SCD(net196),
.SCE(net318),
.SET_B(net308),
.CLK_N(clk),
.Q(net335),
.Q_N(net334)
);

sky130_fd_sc_hd__mux4_1 c424(
.A0(in27),
.A1(net330),
.A2(net335),
.A3(net331),
.S0(net317),
.S1(net329),
.X(net336)
);

sky130_fd_sc_hd__o2111ai_1 c425(
.A1(net220),
.A2(in27),
.B1(net331),
.C1(in29),
.D1(net804),
.Y(net337)
);

sky130_fd_sc_hd__a2111oi_1 c426(
.A1(net332),
.A2(net196),
.B1(net214),
.C1(net334),
.D1(net805),
.Y(net338)
);

sky130_fd_sc_hd__sdfbbn_2 c427(
.D(net329),
.RESET_B(net203),
.SCD(net331),
.SCE(net330),
.SET_B(net220),
.CLK_N(clk),
.Q(net340),
.Q_N(net339)
);

sky130_fd_sc_hd__sdfbbp_1 c428(
.D(net333),
.RESET_B(net209),
.SCD(net318),
.SCE(net334),
.SET_B(net200),
.CLK(clk),
.Q(net342),
.Q_N(net341)
);

sky130_fd_sc_hd__sdfrtp_1 c429(
.D(net340),
.RESET_B(net324),
.SCD(net333),
.SCE(net650),
.CLK(clk),
.Q(net343)
);

sky130_fd_sc_hd__mux4_2 c430(
.A0(net343),
.A1(net315),
.A2(in41),
.A3(net341),
.S0(out1),
.S1(net802),
.X(net344)
);

sky130_fd_sc_hd__mux4_4 c431(
.A0(net196),
.A1(net232),
.A2(net343),
.A3(net333),
.S0(net344),
.S1(net804),
.X(net345)
);

sky130_fd_sc_hd__sdfbbn_1 c432(
.D(net342),
.RESET_B(net331),
.SCD(net209),
.SCE(net343),
.SET_B(net334),
.CLK_N(clk),
.Q(net347),
.Q_N(net346)
);

sky130_fd_sc_hd__mux4_2 c433(
.A0(net316),
.A1(net321),
.A2(net347),
.A3(net339),
.S0(net343),
.S1(net802),
.X(net348)
);

sky130_fd_sc_hd__mux4_4 c434(
.A0(net202),
.A1(net332),
.A2(net340),
.A3(net209),
.S0(net344),
.S1(net650),
.X(net349)
);

sky130_fd_sc_hd__mux4_4 c435(
.A0(net324),
.A1(net232),
.A2(net229),
.A3(net342),
.S0(net321),
.S1(net806),
.X(net350)
);

sky130_fd_sc_hd__mux4_2 c436(
.A0(net81),
.A1(net339),
.A2(net329),
.A3(net315),
.S0(net805),
.S1(out24),
.X(net351)
);

sky130_fd_sc_hd__mux4_1 c437(
.A0(net351),
.A1(net345),
.A2(net333),
.A3(net220),
.S0(net343),
.S1(out24),
.X(net352)
);

sky130_fd_sc_hd__mux4_4 c438(
.A0(net222),
.A1(net332),
.A2(net203),
.A3(net650),
.S0(net800),
.S1(net804),
.X(net353)
);

sky130_fd_sc_hd__mux4_1 c439(
.A0(net348),
.A1(net228),
.A2(net346),
.A3(net232),
.S0(net351),
.S1(net807),
.X(net354)
);

sky130_fd_sc_hd__mux4_4 c440(
.A0(net231),
.A1(net331),
.A2(net332),
.A3(net204),
.S0(in57),
.S1(net676),
.X(net355)
);

sky130_fd_sc_hd__a2111o_1 c441(
.A1(net342),
.A2(in13),
.B1(in52),
.C1(in0),
.D1(net799),
.X(net356)
);

sky130_fd_sc_hd__sdfbbn_2 c442(
.D(net356),
.RESET_B(net237),
.SCD(net331),
.SCE(net214),
.SET_B(in0),
.CLK_N(clk),
.Q(out18),
.Q_N(net357)
);

sky130_fd_sc_hd__or3b_4 c443(
.A(in57),
.B(in52),
.C_N(net249),
.X(net358)
);

sky130_fd_sc_hd__sdfbbp_1 c444(
.D(net358),
.RESET_B(out38),
.SCD(net124),
.SCE(net257),
.SET_B(net785),
.CLK(clk),
.Q(net360),
.Q_N(net359)
);

sky130_fd_sc_hd__or4bb_1 c445(
.A(net245),
.B(net345),
.C_N(net358),
.D_N(in57),
.X(net361)
);

sky130_fd_sc_hd__or4bb_1 c446(
.A(net345),
.B(net734),
.C_N(net750),
.D_N(net758),
.X(net362)
);

sky130_fd_sc_hd__sdfbbn_1 c447(
.D(net360),
.RESET_B(net332),
.SCD(in29),
.SCE(net249),
.SET_B(net808),
.CLK_N(clk),
.Q(net364),
.Q_N(net363)
);

sky130_fd_sc_hd__nor3_2 c448(
.A(net360),
.B(net341),
.C(out24),
.Y(net365)
);

sky130_fd_sc_hd__or4bb_1 c449(
.A(net365),
.B(in0),
.C_N(net749),
.D_N(net783),
.X(net366)
);

sky130_fd_sc_hd__mux4_2 c450(
.A0(net257),
.A1(net359),
.A2(net365),
.A3(net204),
.S0(net346),
.S1(out1),
.X(net367)
);

sky130_fd_sc_hd__mux4_4 c451(
.A0(net124),
.A1(net364),
.A2(net203),
.A3(net97),
.S0(net784),
.S1(net808),
.X(net368)
);

sky130_fd_sc_hd__mux4_2 c452(
.A0(net368),
.A1(in35),
.A2(net363),
.A3(net246),
.S0(net113),
.S1(net684),
.X(net369)
);

sky130_fd_sc_hd__mux4_2 c453(
.A0(net365),
.A1(net359),
.A2(net369),
.A3(net341),
.S0(net212),
.S1(net676),
.X(net370)
);

sky130_fd_sc_hd__mux4_1 c454(
.A0(net347),
.A1(net342),
.A2(net366),
.A3(in41),
.S0(net310),
.S1(out40),
.X(net371)
);

sky130_fd_sc_hd__or4bb_2 c455(
.A(net357),
.B(net113),
.C_N(out40),
.D_N(net785),
.X(net372)
);

sky130_fd_sc_hd__mux4_2 c456(
.A0(in48),
.A1(net346),
.A2(net372),
.A3(net749),
.S0(net758),
.S1(net807),
.X(net373)
);

sky130_fd_sc_hd__a2111o_4 c457(
.A1(net366),
.A2(net371),
.B1(net372),
.C1(net332),
.D1(net713),
.X(net374)
);

sky130_fd_sc_hd__o2111a_2 c458(
.A1(net347),
.A2(net357),
.B1(net684),
.C1(net713),
.D1(out5),
.X(net375)
);

sky130_fd_sc_hd__a2111o_4 c459(
.A1(net371),
.A2(net373),
.B1(net672),
.C1(out1),
.D1(net807),
.X(net376)
);

sky130_fd_sc_hd__mux4_2 c460(
.A0(net375),
.A1(in2),
.A2(net363),
.A3(net372),
.S0(net376),
.S1(net672),
.X(net377)
);

sky130_fd_sc_hd__o2111ai_1 c461(
.A1(net242),
.A2(net377),
.B1(net376),
.C1(net368),
.D1(net375),
.Y(net378)
);

sky130_fd_sc_hd__mux4_1 c462(
.A0(net315),
.A1(net377),
.A2(out31),
.A3(net12),
.S0(net284),
.S1(net807),
.X(out4)
);

sky130_fd_sc_hd__mux4_4 c463(
.A0(net12),
.A1(out18),
.A2(net209),
.A3(net378),
.S0(net792),
.S1(net800),
.X(net379)
);

sky130_fd_sc_hd__mux4_4 c464(
.A0(out4),
.A1(in4),
.A2(net372),
.A3(net778),
.S0(net795),
.S1(net808),
.X(net380)
);

sky130_fd_sc_hd__mux4_2 c465(
.A0(net377),
.A1(net330),
.A2(net331),
.A3(net372),
.S0(net738),
.S1(net787),
.X(net381)
);

sky130_fd_sc_hd__mux4_4 c466(
.A0(net281),
.A1(in31),
.A2(net97),
.A3(net378),
.S0(net808),
.S1(net810),
.X(net382)
);

sky130_fd_sc_hd__mux4_4 c467(
.A0(net369),
.A1(net377),
.A2(net793),
.A3(net795),
.S0(net799),
.S1(out24),
.X(net383)
);

sky130_fd_sc_hd__mux4_4 c468(
.A0(net369),
.A1(out4),
.A2(net738),
.A3(net793),
.S0(net807),
.S1(net810),
.X(net384)
);

sky130_fd_sc_hd__mux4_2 c469(
.A0(net330),
.A1(net329),
.A2(out49),
.A3(net793),
.S0(out39),
.S1(net809),
.X(net385)
);

sky130_fd_sc_hd__mux4_4 c470(
.A0(out31),
.A1(net77),
.A2(out42),
.A3(out24),
.S0(out39),
.S1(net810),
.X(net386)
);

sky130_fd_sc_hd__mux4_4 c471(
.A0(net378),
.A1(out42),
.A2(net801),
.A3(net807),
.S0(out39),
.S1(net809),
.X(net387)
);

sky130_fd_sc_hd__mux4_2 c472(
.A0(net330),
.A1(out4),
.A2(net738),
.A3(net788),
.S0(net808),
.S1(out39),
.X(net388)
);

sky130_fd_sc_hd__mux4_1 c473(
.A0(net331),
.A1(net369),
.A2(net18),
.A3(net738),
.S0(net792),
.S1(net799),
.X(net389)
);

sky130_fd_sc_hd__mux4_1 c474(
.A0(out38),
.A1(net19),
.A2(net738),
.A3(out7),
.S0(out39),
.S1(net812),
.X(net390)
);

sky130_fd_sc_hd__mux4_2 c475(
.A0(out38),
.A1(out49),
.A2(out1),
.A3(net785),
.S0(out39),
.S1(net809),
.X(net391)
);

sky130_fd_sc_hd__mux4_1 c476(
.A0(net329),
.A1(net391),
.A2(net281),
.A3(net386),
.S0(net787),
.S1(net810),
.X(net392)
);

sky130_fd_sc_hd__mux4_1 c477(
.A0(net7),
.A1(net391),
.A2(net12),
.A3(out42),
.S0(net812),
.S1(out9),
.X(net393)
);

sky130_fd_sc_hd__mux4_4 c478(
.A0(net391),
.A1(net393),
.A2(in48),
.A3(net801),
.S0(net811),
.S1(out9),
.X(net394)
);

sky130_fd_sc_hd__mux4_4 c479(
.A0(net393),
.A1(out4),
.A2(net330),
.A3(net799),
.S0(net807),
.S1(net812),
.X(net395)
);

sky130_fd_sc_hd__mux4_4 c480(
.A0(net390),
.A1(net391),
.A2(net245),
.A3(net281),
.S0(out39),
.S1(net811),
.X(net396)
);

sky130_fd_sc_hd__mux4_2 c481(
.A0(net396),
.A1(in46),
.A2(net391),
.A3(out31),
.S0(net784),
.S1(net795),
.X(net397)
);

sky130_fd_sc_hd__mux4_2 c482(
.A0(net397),
.A1(in46),
.A2(out31),
.A3(net738),
.S0(out9),
.S1(net813),
.X(net398)
);

sky130_fd_sc_hd__mux4_1 c483(
.A0(net391),
.A1(net396),
.A2(net397),
.A3(out49),
.S0(out9),
.S1(net813),
.X(net399)
);

sky130_fd_sc_hd__mux4_2 c484(
.A0(out18),
.A1(net300),
.A2(net771),
.A3(net796),
.S0(net798),
.S1(out24),
.X(net400)
);

sky130_fd_sc_hd__mux4_2 c485(
.A0(in48),
.A1(net300),
.A2(out32),
.A3(out25),
.S0(net34),
.S1(out39),
.X(net401)
);

sky130_fd_sc_hd__mux4_2 c486(
.A0(net377),
.A1(net329),
.A2(net295),
.A3(out12),
.S0(net768),
.S1(out39),
.X(net402)
);

sky130_fd_sc_hd__mux4_1 c487(
.A0(net401),
.A1(net339),
.A2(net764),
.A3(net768),
.S0(net769),
.S1(net770),
.X(net403)
);

sky130_fd_sc_hd__mux4_4 c488(
.A0(net119),
.A1(net340),
.A2(in61),
.A3(net403),
.S0(net34),
.S1(net787),
.X(net404)
);

sky130_fd_sc_hd__mux4_4 c489(
.A0(net403),
.A1(net18),
.A2(net113),
.A3(out31),
.S0(net401),
.S1(net300),
.X(net405)
);

sky130_fd_sc_hd__mux4_2 c490(
.A0(net401),
.A1(net296),
.A2(net300),
.A3(net403),
.S0(net698),
.S1(net735),
.X(net406)
);

sky130_fd_sc_hd__mux4_4 c491(
.A0(in52),
.A1(out31),
.A2(net401),
.A3(out30),
.S0(net762),
.S1(out13),
.X(out8)
);

sky130_fd_sc_hd__mux4_2 c492(
.A0(net400),
.A1(net403),
.A2(out16),
.A3(net104),
.S0(out30),
.S1(out39),
.X(net407)
);

sky130_fd_sc_hd__mux4_4 c493(
.A0(net403),
.A1(out29),
.A2(net735),
.A3(out15),
.S0(net768),
.S1(net815),
.X(net408)
);

sky130_fd_sc_hd__mux4_1 c494(
.A0(net302),
.A1(net403),
.A2(net401),
.A3(net814),
.S0(net815),
.S1(out10),
.X(net409)
);

sky130_fd_sc_hd__mux4_4 c495(
.A0(out25),
.A1(out8),
.A2(out38),
.A3(net735),
.S0(net798),
.S1(net816),
.X(net410)
);

sky130_fd_sc_hd__mux4_4 c496(
.A0(net303),
.A1(net209),
.A2(out29),
.A3(net403),
.S0(out30),
.S1(net763),
.X(net411)
);

sky130_fd_sc_hd__mux4_1 c497(
.A0(net329),
.A1(out8),
.A2(net403),
.A3(out15),
.S0(net796),
.S1(net815),
.X(net412)
);

sky130_fd_sc_hd__mux4_4 c498(
.A0(net340),
.A1(out8),
.A2(out49),
.A3(net770),
.S0(net798),
.S1(net818),
.X(net413)
);

sky130_fd_sc_hd__mux4_1 c499(
.A0(out32),
.A1(net403),
.A2(net768),
.A3(net771),
.S0(net787),
.S1(net819),
.X(net414)
);

sky130_fd_sc_hd__mux4_1 c500(
.A0(net115),
.A1(net213),
.A2(out25),
.A3(out12),
.S0(net735),
.S1(net815),
.X(net415)
);

sky130_fd_sc_hd__mux4_2 c501(
.A0(out32),
.A1(net735),
.A2(net787),
.A3(out13),
.S0(net819),
.S1(net821),
.X(out41)
);

sky130_fd_sc_hd__mux4_4 c502(
.A0(net34),
.A1(net115),
.A2(net735),
.A3(net770),
.S0(net814),
.S1(net820),
.X(out34)
);

sky130_fd_sc_hd__mux4_4 c503(
.A0(net372),
.A1(out34),
.A2(net401),
.A3(out41),
.S0(out40),
.S1(net820),
.X(out23)
);

sky130_fd_sc_hd__mux4_4 c504(
.A0(out34),
.A1(out23),
.A2(out41),
.A3(out8),
.S0(out49),
.S1(net818),
.X(net416)
);

sky130_fd_sc_hd__mux4_4 c505(
.A0(net104),
.A1(out34),
.A2(out23),
.A3(out29),
.S0(net403),
.S1(net725),
.X(net417)
);

sky130_fd_sc_hd__or3b_4 c528(
.A(net207),
.B(net312),
.C_N(net320),
.X(net418)
);

sky130_fd_sc_hd__nor3b_2 c529(
.A(net72),
.B(net320),
.C_N(in0),
.Y(net419)
);

sky130_fd_sc_hd__and3_4 c530(
.A(net328),
.B(net201),
.C(in0),
.X(net420)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c531(
.A(net737),
.X(out14)
);

sky130_fd_sc_hd__a2111oi_0 c532(
.A1(net201),
.A2(net328),
.B1(net203),
.C1(net321),
.D1(net803),
.Y(net421)
);

sky130_fd_sc_hd__dlygate4sd3_1 c533(
.A(net737),
.X(net422)
);

sky130_fd_sc_hd__buf_16 c534(
.A(net706),
.X(net423)
);

sky130_fd_sc_hd__inv_6 c535(
.A(net737),
.Y(net424)
);

sky130_fd_sc_hd__nor3b_1 c536(
.A(net424),
.B(net422),
.C_N(net423),
.Y(out2)
);

sky130_fd_sc_hd__inv_1 c537(
.A(net706),
.Y(net425)
);

sky130_fd_sc_hd__sdfrtp_2 c538(
.D(net423),
.RESET_B(net312),
.SCD(net328),
.SCE(net419),
.CLK(clk),
.Q(net426)
);

sky130_fd_sc_hd__a2111o_4 c539(
.A1(net208),
.A2(net425),
.B1(net420),
.C1(net422),
.D1(in0),
.X(net427)
);

sky130_fd_sc_hd__sdfbbn_2 c540(
.D(net419),
.RESET_B(net425),
.SCD(net310),
.SCE(net217),
.SET_B(net426),
.CLK_N(clk),
.Q(net429),
.Q_N(net428)
);

sky130_fd_sc_hd__clkbuf_2 c541(
.A(net737),
.X(net430)
);

sky130_fd_sc_hd__or3_1 c542(
.A(net429),
.B(net430),
.C(net426),
.X(net431)
);

sky130_fd_sc_hd__mux4_4 c543(
.A0(net426),
.A1(net428),
.A2(net425),
.A3(out14),
.S0(net207),
.S1(net418),
.X(net432)
);

sky130_fd_sc_hd__mux4_2 c544(
.A0(net422),
.A1(out2),
.A2(net425),
.A3(net321),
.S0(net318),
.S1(net803),
.X(net433)
);

sky130_fd_sc_hd__mux4_2 c545(
.A0(net423),
.A1(net426),
.A2(net321),
.A3(net419),
.S0(in4),
.S1(net424),
.X(net434)
);

sky130_fd_sc_hd__mux4_4 c546(
.A0(net217),
.A1(net424),
.A2(net433),
.A3(net723),
.S0(net726),
.S1(net822),
.X(net435)
);

sky130_fd_sc_hd__mux4_4 c547(
.A0(net433),
.A1(net431),
.A2(net424),
.A3(net425),
.S0(net321),
.S1(net822),
.X(net436)
);

sky130_fd_sc_hd__mux4_4 c548(
.A0(net433),
.A1(net428),
.A2(net419),
.A3(net723),
.S0(net730),
.S1(net823),
.X(net437)
);

sky130_fd_sc_hd__mux4_2 c549(
.A0(in2),
.A1(net318),
.A2(net422),
.A3(net420),
.S0(net730),
.S1(net737),
.X(net438)
);

sky130_fd_sc_hd__a2111o_4 c550(
.A1(net318),
.A2(net335),
.B1(net344),
.C1(out24),
.D1(net823),
.X(net439)
);

sky130_fd_sc_hd__or4bb_4 c551(
.A(in29),
.B(net318),
.C_N(in37),
.D_N(net76),
.X(net440)
);

sky130_fd_sc_hd__a2111oi_2 c552(
.A1(net439),
.A2(net318),
.B1(net228),
.C1(net440),
.D1(net805),
.Y(net441)
);

sky130_fd_sc_hd__nand3_2 c553(
.A(net335),
.B(in37),
.C(net823),
.Y(net442)
);

sky130_fd_sc_hd__o2111ai_4 c554(
.A1(net442),
.A2(net335),
.B1(in2),
.C1(net726),
.D1(out24),
.Y(net443)
);

sky130_fd_sc_hd__o2111ai_1 c555(
.A1(net237),
.A2(net441),
.B1(net334),
.C1(net726),
.D1(net804),
.Y(net444)
);

sky130_fd_sc_hd__or4bb_1 c556(
.A(net443),
.B(in0),
.C_N(net685),
.D_N(net757),
.X(net445)
);

sky130_fd_sc_hd__or3_4 c557(
.A(net328),
.B(net442),
.C(net806),
.X(net446)
);

sky130_fd_sc_hd__or4bb_1 c558(
.A(net321),
.B(net335),
.C_N(net222),
.D_N(net822),
.X(net447)
);

sky130_fd_sc_hd__sdfrtp_4 c559(
.D(net439),
.RESET_B(net441),
.SCD(net237),
.SCE(net442),
.CLK(clk),
.Q(out11)
);

sky130_fd_sc_hd__mux4_1 c560(
.A0(net429),
.A1(net228),
.A2(in35),
.A3(net650),
.S0(net805),
.S1(net806),
.X(net448)
);

sky130_fd_sc_hd__a2111oi_4 c561(
.A1(net446),
.A2(net228),
.B1(in0),
.C1(net447),
.D1(net757),
.Y(net449)
);

sky130_fd_sc_hd__a2111o_1 c562(
.A1(net445),
.A2(net428),
.B1(net439),
.C1(net76),
.D1(net804),
.X(net450)
);

sky130_fd_sc_hd__sdfbbp_1 c563(
.D(out11),
.RESET_B(net447),
.SCD(net445),
.SCE(net318),
.SET_B(net685),
.CLK(clk),
.Q(net452),
.Q_N(net451)
);

sky130_fd_sc_hd__o2111ai_4 c564(
.A1(net429),
.A2(net443),
.B1(net452),
.C1(net318),
.D1(net448),
.Y(net453)
);

sky130_fd_sc_hd__sdfbbn_1 c565(
.D(net453),
.RESET_B(net421),
.SCD(net439),
.SCE(net447),
.SET_B(net228),
.CLK_N(clk),
.Q(net455),
.Q_N(net454)
);

sky130_fd_sc_hd__a2111o_2 c566(
.A1(net222),
.A2(net454),
.B1(net757),
.C1(net802),
.D1(net805),
.X(out17)
);

sky130_fd_sc_hd__mux4_1 c567(
.A0(net441),
.A1(net452),
.A2(net454),
.A3(net439),
.S0(out11),
.S1(net447),
.X(net456)
);

sky130_fd_sc_hd__or4bb_1 c568(
.A(net447),
.B(net455),
.C_N(out17),
.D_N(net451),
.X(net457)
);

sky130_fd_sc_hd__mux4_4 c569(
.A0(net450),
.A1(net447),
.A2(net310),
.A3(net685),
.S0(net726),
.S1(net806),
.X(net458)
);

sky130_fd_sc_hd__mux4_1 c570(
.A0(net447),
.A1(net454),
.A2(net451),
.A3(net453),
.S0(net685),
.S1(net825),
.X(net459)
);

sky130_fd_sc_hd__mux4_1 c571(
.A0(net440),
.A1(net231),
.A2(net446),
.A3(net726),
.S0(net805),
.S1(out21),
.X(net460)
);

sky130_fd_sc_hd__mux4_4 c572(
.A0(net376),
.A1(out2),
.A2(in29),
.A3(net249),
.S0(net310),
.S1(net822),
.X(net461)
);

sky130_fd_sc_hd__mux4_4 c573(
.A0(net246),
.A1(net440),
.A2(net422),
.A3(in61),
.S0(net448),
.S1(net368),
.X(net462)
);

sky130_fd_sc_hd__mux4_4 c574(
.A0(net76),
.A1(net373),
.A2(net462),
.A3(net369),
.S0(net378),
.S1(net372),
.X(net463)
);

sky130_fd_sc_hd__mux4_1 c575(
.A0(net368),
.A1(net203),
.A2(out5),
.A3(net778),
.S0(net806),
.S1(net826),
.X(net464)
);

sky130_fd_sc_hd__mux4_2 c576(
.A0(net364),
.A1(net104),
.A2(net310),
.A3(out2),
.S0(net249),
.S1(net783),
.X(net465)
);

sky130_fd_sc_hd__mux4_2 c577(
.A0(net440),
.A1(net462),
.A2(net376),
.A3(in2),
.S0(net465),
.S1(net122),
.X(net466)
);

sky130_fd_sc_hd__mux4_4 c578(
.A0(net373),
.A1(net104),
.A2(net726),
.A3(net806),
.S0(out21),
.S1(net828),
.X(net467)
);

sky130_fd_sc_hd__mux4_2 c579(
.A0(net310),
.A1(net373),
.A2(net465),
.A3(net97),
.S0(net462),
.S1(net376),
.X(net468)
);

sky130_fd_sc_hd__mux4_1 c580(
.A0(net452),
.A1(net372),
.A2(net104),
.A3(net461),
.S0(net806),
.S1(net828),
.X(net469)
);

sky130_fd_sc_hd__mux4_1 c581(
.A0(net310),
.A1(net372),
.A2(net462),
.A3(net465),
.S0(net824),
.S1(net829),
.X(net470)
);

sky130_fd_sc_hd__mux4_2 c582(
.A0(net373),
.A1(net465),
.A2(in35),
.A3(net822),
.S0(net826),
.S1(net830),
.X(net471)
);

sky130_fd_sc_hd__mux4_4 c583(
.A0(net464),
.A1(net373),
.A2(net471),
.A3(net698),
.S0(net713),
.S1(net822),
.X(net472)
);

sky130_fd_sc_hd__mux4_1 c584(
.A0(net471),
.A1(net213),
.A2(net364),
.A3(net72),
.S0(net373),
.S1(net830),
.X(net473)
);

sky130_fd_sc_hd__mux4_4 c585(
.A0(net373),
.A1(net461),
.A2(in41),
.A3(net715),
.S0(net758),
.S1(net830),
.X(net474)
);

sky130_fd_sc_hd__mux4_1 c586(
.A0(out14),
.A1(net246),
.A2(net825),
.A3(out21),
.S0(net830),
.S1(net831),
.X(net475)
);

sky130_fd_sc_hd__mux4_4 c587(
.A0(net465),
.A1(net461),
.A2(net203),
.A3(net475),
.S0(net469),
.S1(net462),
.X(net476)
);

sky130_fd_sc_hd__mux4_2 c588(
.A0(net249),
.A1(net474),
.A2(net475),
.A3(net825),
.S0(net829),
.S1(net831),
.X(net477)
);

sky130_fd_sc_hd__mux4_1 c589(
.A0(out18),
.A1(net76),
.A2(net310),
.A3(net465),
.S0(net475),
.S1(net737),
.X(net478)
);

sky130_fd_sc_hd__mux4_4 c590(
.A0(net475),
.A1(net378),
.A2(out1),
.A3(out24),
.S0(net829),
.S1(net830),
.X(net479)
);

sky130_fd_sc_hd__mux4_2 c591(
.A0(net475),
.A1(net469),
.A2(net715),
.A3(net724),
.S0(net758),
.S1(out24),
.X(net480)
);

sky130_fd_sc_hd__mux4_4 c592(
.A0(net115),
.A1(net684),
.A2(net717),
.A3(net724),
.S0(net737),
.S1(out21),
.X(net481)
);

sky130_fd_sc_hd__mux4_1 c593(
.A0(net469),
.A1(net475),
.A2(net481),
.A3(net465),
.S0(net717),
.S1(net724),
.X(net482)
);

sky130_fd_sc_hd__mux4_2 c594(
.A0(net19),
.A1(net448),
.A2(out14),
.A3(out2),
.S0(in4),
.S1(net77),
.X(net483)
);

sky130_fd_sc_hd__mux4_1 c595(
.A0(net467),
.A1(net372),
.A2(net249),
.A3(out7),
.S0(net789),
.S1(out9),
.X(net484)
);

sky130_fd_sc_hd__mux4_4 c596(
.A0(net448),
.A1(out2),
.A2(net789),
.A3(out24),
.S0(out21),
.S1(net827),
.X(net485)
);

sky130_fd_sc_hd__mux4_2 c597(
.A0(net19),
.A1(out14),
.A2(net483),
.A3(net717),
.S0(net788),
.S1(net814),
.X(net486)
);

sky130_fd_sc_hd__mux4_1 c598(
.A0(net203),
.A1(net19),
.A2(net684),
.A3(out49),
.S0(net783),
.S1(net831),
.X(net487)
);

sky130_fd_sc_hd__mux4_4 c599(
.A0(net461),
.A1(net394),
.A2(net19),
.A3(out4),
.S0(net77),
.S1(net814),
.X(net488)
);

sky130_fd_sc_hd__mux4_2 c600(
.A0(net486),
.A1(in46),
.A2(net372),
.A3(net454),
.S0(net721),
.S1(net831),
.X(net489)
);

sky130_fd_sc_hd__mux4_1 c601(
.A0(net448),
.A1(net344),
.A2(out2),
.A3(out14),
.S0(net212),
.S1(net831),
.X(net490)
);

sky130_fd_sc_hd__mux4_4 c602(
.A0(net484),
.A1(net19),
.A2(net249),
.A3(net481),
.S0(net212),
.S1(net826),
.X(net491)
);

sky130_fd_sc_hd__mux4_2 c603(
.A0(net487),
.A1(net481),
.A2(in4),
.A3(net721),
.S0(net731),
.S1(out9),
.X(net492)
);

sky130_fd_sc_hd__mux4_1 c604(
.A0(net490),
.A1(net77),
.A2(net467),
.A3(net483),
.S0(net731),
.S1(net789),
.X(net493)
);

sky130_fd_sc_hd__mux4_2 c605(
.A0(net493),
.A1(net394),
.A2(net284),
.A3(net487),
.S0(net77),
.S1(net721),
.X(net494)
);

sky130_fd_sc_hd__mux4_2 c606(
.A0(net493),
.A1(net104),
.A2(net492),
.A3(net487),
.S0(net372),
.S1(out24),
.X(net495)
);

sky130_fd_sc_hd__mux4_1 c607(
.A0(net485),
.A1(net492),
.A2(net237),
.A3(net378),
.S0(net789),
.S1(net833),
.X(net496)
);

sky130_fd_sc_hd__mux4_2 c608(
.A0(net394),
.A1(net493),
.A2(net683),
.A3(net783),
.S0(net831),
.S1(net833),
.X(net497)
);

sky130_fd_sc_hd__mux4_2 c609(
.A0(in29),
.A1(net487),
.A2(net788),
.A3(out39),
.S0(net833),
.S1(net835),
.X(net498)
);

sky130_fd_sc_hd__mux4_2 c610(
.A0(net498),
.A1(net483),
.A2(net19),
.A3(net683),
.S0(net833),
.S1(net835),
.X(net499)
);

sky130_fd_sc_hd__mux4_1 c611(
.A0(net113),
.A1(net97),
.A2(net498),
.A3(net481),
.S0(net731),
.S1(out1),
.X(net500)
);

sky130_fd_sc_hd__mux4_2 c612(
.A0(net499),
.A1(net249),
.A2(net498),
.A3(net490),
.S0(net378),
.S1(net835),
.X(net501)
);

sky130_fd_sc_hd__mux4_1 c613(
.A0(net378),
.A1(net487),
.A2(net394),
.A3(net483),
.S0(net834),
.S1(net836),
.X(net502)
);

sky130_fd_sc_hd__mux4_1 c614(
.A0(net492),
.A1(net499),
.A2(net490),
.A3(net682),
.S0(net831),
.S1(net835),
.X(net503)
);

sky130_fd_sc_hd__mux4_4 c615(
.A0(net498),
.A1(net500),
.A2(net487),
.A3(net490),
.S0(net682),
.S1(net837),
.X(net504)
);

sky130_fd_sc_hd__mux4_2 c616(
.A0(net18),
.A1(net249),
.A2(net821),
.A3(net827),
.S0(out19),
.S1(net838),
.X(net505)
);

sky130_fd_sc_hd__mux4_2 c617(
.A0(net481),
.A1(net505),
.A2(net771),
.A3(net788),
.S0(out13),
.S1(net839),
.X(net506)
);

sky130_fd_sc_hd__mux4_4 c618(
.A0(net34),
.A1(out2),
.A2(out24),
.A3(out39),
.S0(net827),
.S1(net833),
.X(net507)
);

sky130_fd_sc_hd__mux4_2 c619(
.A0(net506),
.A1(net18),
.A2(net357),
.A3(out16),
.S0(out13),
.S1(net834),
.X(net508)
);

sky130_fd_sc_hd__mux4_1 c620(
.A0(net34),
.A1(out8),
.A2(net769),
.A3(net815),
.S0(net826),
.S1(net831),
.X(net509)
);

sky130_fd_sc_hd__mux4_1 c621(
.A0(net508),
.A1(net372),
.A2(out14),
.A3(out15),
.S0(net788),
.S1(net839),
.X(net510)
);

sky130_fd_sc_hd__mux4_4 c622(
.A0(net300),
.A1(net506),
.A2(out15),
.A3(out9),
.S0(net816),
.S1(net833),
.X(net511)
);

sky130_fd_sc_hd__mux4_1 c623(
.A0(net506),
.A1(net508),
.A2(out2),
.A3(net769),
.S0(out7),
.S1(out10),
.X(net512)
);

sky130_fd_sc_hd__mux4_1 c624(
.A0(net511),
.A1(net481),
.A2(in61),
.A3(out10),
.S0(net827),
.S1(net838),
.X(net513)
);

sky130_fd_sc_hd__mux4_1 c625(
.A0(net512),
.A1(net34),
.A2(net213),
.A3(out11),
.S0(net820),
.S1(out3),
.X(net514)
);

sky130_fd_sc_hd__mux4_2 c626(
.A0(net104),
.A1(net122),
.A2(net483),
.A3(net34),
.S0(net510),
.S1(net827),
.X(net515)
);

sky130_fd_sc_hd__mux4_4 c627(
.A0(net481),
.A1(net113),
.A2(out14),
.A3(net698),
.S0(net716),
.S1(out10),
.X(net516)
);

sky130_fd_sc_hd__mux4_2 c628(
.A0(net508),
.A1(out16),
.A2(in61),
.A3(net762),
.S0(net771),
.S1(net788),
.X(out20)
);

sky130_fd_sc_hd__mux4_1 c629(
.A0(net455),
.A1(net507),
.A2(net483),
.A3(out14),
.S0(out13),
.S1(net836),
.X(net517)
);

sky130_fd_sc_hd__mux4_2 c630(
.A0(net516),
.A1(net515),
.A2(net517),
.A3(net212),
.S0(net762),
.S1(net834),
.X(net518)
);

sky130_fd_sc_hd__mux4_1 c631(
.A0(net455),
.A1(in13),
.A2(net698),
.A3(out1),
.S0(net833),
.S1(net834),
.X(out6)
);

sky130_fd_sc_hd__mux4_2 c632(
.A0(in41),
.A1(out6),
.A2(net510),
.A3(net814),
.S0(net817),
.S1(out19),
.X(out0)
);

sky130_fd_sc_hd__mux4_1 c633(
.A0(net513),
.A1(net517),
.A2(out0),
.A3(net300),
.S0(net508),
.S1(net722),
.X(net519)
);

sky130_fd_sc_hd__mux4_2 c634(
.A0(net517),
.A1(out0),
.A2(net510),
.A3(net716),
.S0(net722),
.S1(net834),
.X(net520)
);

sky130_fd_sc_hd__mux4_4 c635(
.A0(net213),
.A1(in61),
.A2(net717),
.A3(out15),
.S0(net798),
.S1(net834),
.X(net521)
);

sky130_fd_sc_hd__mux4_2 c636(
.A0(net521),
.A1(out17),
.A2(out0),
.A3(net762),
.S0(net814),
.S1(net836),
.X(net522)
);

sky130_fd_sc_hd__mux4_2 c637(
.A0(net514),
.A1(net284),
.A2(net515),
.A3(net510),
.S0(net517),
.S1(net722),
.X(net523)
);

sky130_fd_sc_hd__inv_12 c660(
.A(net696),
.Y(net524)
);

sky130_fd_sc_hd__inv_4 c661(
.A(net696),
.Y(net525)
);

sky130_fd_sc_hd__nor3b_4 c662(
.A(net431),
.B(net525),
.C_N(net320),
.Y(net526)
);

sky130_fd_sc_hd__mux4_4 c663(
.A0(net81),
.A1(net422),
.A2(net77),
.A3(net328),
.S0(net525),
.S1(net418),
.X(net527)
);

sky130_fd_sc_hd__buf_8 c664(
.A(net719),
.X(net528)
);

sky130_fd_sc_hd__nor3_1 c665(
.A(net312),
.B(net424),
.C(net528),
.Y(net529)
);

sky130_fd_sc_hd__and3_1 c666(
.A(net528),
.B(net525),
.C(net529),
.X(net530)
);

sky130_fd_sc_hd__nor3b_4 c667(
.A(net320),
.B(net312),
.C_N(net823),
.Y(net531)
);

sky130_fd_sc_hd__mux4_1 c668(
.A0(net529),
.A1(net214),
.A2(net525),
.A3(net320),
.S0(net528),
.S1(net723),
.X(net532)
);

sky130_fd_sc_hd__buf_2 c669(
.A(net719),
.X(net533)
);

sky130_fd_sc_hd__mux4_1 c670(
.A0(net532),
.A1(net312),
.A2(net533),
.A3(net425),
.S0(net422),
.S1(net525),
.X(net534)
);

sky130_fd_sc_hd__or3_2 c671(
.A(net533),
.B(net312),
.C(net730),
.X(net535)
);

sky130_fd_sc_hd__mux4_1 c672(
.A0(net530),
.A1(net531),
.A2(net533),
.A3(net525),
.S0(net528),
.S1(net841),
.X(net536)
);

sky130_fd_sc_hd__o2111a_2 c673(
.A1(net532),
.A2(net528),
.B1(net535),
.C1(net533),
.D1(net525),
.X(net537)
);

sky130_fd_sc_hd__or4bb_2 c674(
.A(net217),
.B(net533),
.C_N(net528),
.D_N(net728),
.X(net538)
);

sky130_fd_sc_hd__mux4_1 c675(
.A0(net430),
.A1(net530),
.A2(in0),
.A3(net533),
.S0(net431),
.S1(net532),
.X(net539)
);

sky130_fd_sc_hd__mux4_2 c676(
.A0(net419),
.A1(net533),
.A2(net525),
.A3(net728),
.S0(net742),
.S1(net841),
.X(net540)
);

sky130_fd_sc_hd__clkbuf_2 c677(
.A(net719),
.X(net541)
);

sky130_fd_sc_hd__a2111oi_4 c678(
.A1(net528),
.A2(net696),
.B1(net728),
.C1(net742),
.D1(net841),
.Y(net542)
);

sky130_fd_sc_hd__nand3b_4 c679(
.A_N(net529),
.B(net535),
.C(net542),
.Y(net543)
);

sky130_fd_sc_hd__inv_8 c680(
.A(net719),
.Y(net544)
);

sky130_fd_sc_hd__mux4_4 c681(
.A0(net544),
.A1(net531),
.A2(net524),
.A3(net525),
.S0(net528),
.S1(net742),
.X(net545)
);

sky130_fd_sc_hd__o2111a_4 c682(
.A1(net447),
.A2(net525),
.B1(in0),
.C1(net696),
.D1(net778),
.X(net546)
);

sky130_fd_sc_hd__or4bb_4 c683(
.A(net525),
.B(net422),
.C_N(net700),
.D_N(net841),
.X(net547)
);

sky130_fd_sc_hd__or4bb_2 c684(
.A(net524),
.B(in41),
.C_N(net547),
.D_N(net528),
.X(net548)
);

sky130_fd_sc_hd__mux4_2 c685(
.A0(net421),
.A1(net542),
.A2(net443),
.A3(net328),
.S0(in31),
.S1(net842),
.X(net549)
);

sky130_fd_sc_hd__o2111ai_4 c686(
.A1(net344),
.A2(net441),
.B1(net422),
.C1(net542),
.D1(net823),
.Y(net550)
);

sky130_fd_sc_hd__mux4_1 c687(
.A0(net530),
.A1(net525),
.A2(net528),
.A3(net443),
.S0(net228),
.S1(net748),
.X(net551)
);

sky130_fd_sc_hd__o2111ai_2 c688(
.A1(in2),
.A2(net528),
.B1(net542),
.C1(net748),
.D1(net825),
.Y(net552)
);

sky130_fd_sc_hd__a2111oi_0 c689(
.A1(net543),
.A2(net443),
.B1(net344),
.C1(net447),
.D1(net742),
.Y(net553)
);

sky130_fd_sc_hd__o2111ai_1 c690(
.A1(net551),
.A2(net422),
.B1(in0),
.C1(net547),
.D1(net748),
.Y(net554)
);

sky130_fd_sc_hd__sdfbbn_2 c691(
.D(net526),
.RESET_B(net554),
.SCD(in23),
.SCE(net823),
.SET_B(net825),
.CLK_N(clk),
.Q(net556),
.Q_N(net555)
);

sky130_fd_sc_hd__mux4_1 c692(
.A0(net548),
.A1(net555),
.A2(net525),
.A3(net422),
.S0(net344),
.S1(net653),
.X(net557)
);

sky130_fd_sc_hd__or4bb_2 c693(
.A(net525),
.B(net551),
.C_N(net78),
.D_N(net528),
.X(net558)
);

sky130_fd_sc_hd__mux4_2 c694(
.A0(net552),
.A1(net344),
.A2(net441),
.A3(net214),
.S0(net554),
.S1(net547),
.X(net559)
);

sky130_fd_sc_hd__a2111oi_2 c695(
.A1(net548),
.A2(net528),
.B1(net344),
.C1(net653),
.D1(net742),
.Y(net560)
);

sky130_fd_sc_hd__mux4_1 c696(
.A0(net535),
.A1(net528),
.A2(net525),
.A3(net344),
.S0(net551),
.S1(net753),
.X(net561)
);

sky130_fd_sc_hd__o2111ai_4 c697(
.A1(net552),
.A2(net422),
.B1(net560),
.C1(net742),
.D1(net841),
.Y(net562)
);

sky130_fd_sc_hd__mux4_1 c698(
.A0(net556),
.A1(net561),
.A2(net81),
.A3(net447),
.S0(in35),
.S1(net741),
.X(net563)
);

sky130_fd_sc_hd__o2111ai_2 c699(
.A1(net443),
.A2(net441),
.B1(net555),
.C1(net228),
.D1(net843),
.Y(net564)
);

sky130_fd_sc_hd__a2111oi_1 c700(
.A1(net562),
.A2(net447),
.B1(net560),
.C1(net653),
.D1(net843),
.Y(net565)
);

sky130_fd_sc_hd__mux4_1 c701(
.A0(net558),
.A1(net562),
.A2(net552),
.A3(net729),
.S0(net842),
.S1(net843),
.X(net566)
);

sky130_fd_sc_hd__mux4_1 c702(
.A0(net228),
.A1(net447),
.A2(net562),
.A3(net524),
.S0(net729),
.S1(net844),
.X(net567)
);

sky130_fd_sc_hd__mux4_1 c703(
.A0(net560),
.A1(in37),
.A2(net729),
.A3(net754),
.S0(net844),
.S1(net845),
.X(net568)
);

sky130_fd_sc_hd__mux4_2 c704(
.A0(net554),
.A1(net557),
.A2(net328),
.A3(net556),
.S0(net344),
.S1(net824),
.X(net569)
);

sky130_fd_sc_hd__mux4_1 c705(
.A0(net558),
.A1(net203),
.A2(net122),
.A3(in37),
.S0(net344),
.S1(net754),
.X(net570)
);

sky130_fd_sc_hd__mux4_2 c706(
.A0(net424),
.A1(net203),
.A2(in13),
.A3(net824),
.S0(net841),
.S1(net846),
.X(net571)
);

sky130_fd_sc_hd__mux4_4 c707(
.A0(net547),
.A1(net344),
.A2(net474),
.A3(net557),
.S0(net720),
.S1(net841),
.X(net572)
);

sky130_fd_sc_hd__mux4_2 c708(
.A0(net561),
.A1(net215),
.A2(net528),
.A3(net422),
.S0(net832),
.S1(net847),
.X(net573)
);

sky130_fd_sc_hd__mux4_4 c709(
.A0(net474),
.A1(net376),
.A2(in0),
.A3(net841),
.S0(net848),
.S1(net849),
.X(net574)
);

sky130_fd_sc_hd__mux4_4 c710(
.A0(net557),
.A1(net568),
.A2(net474),
.A3(net215),
.S0(net555),
.S1(net849),
.X(net575)
);

sky130_fd_sc_hd__mux4_4 c711(
.A0(net424),
.A1(net77),
.A2(net328),
.A3(net653),
.S0(net832),
.S1(net849),
.X(net576)
);

sky130_fd_sc_hd__mux4_4 c712(
.A0(net376),
.A1(net749),
.A2(net832),
.A3(net841),
.S0(net842),
.S1(net845),
.X(net577)
);

sky130_fd_sc_hd__mux4_4 c713(
.A0(net376),
.A1(net558),
.A2(in2),
.A3(in46),
.S0(net824),
.S1(net851),
.X(net578)
);

sky130_fd_sc_hd__mux4_4 c714(
.A0(net571),
.A1(net576),
.A2(net344),
.A3(net541),
.S0(net845),
.S1(net849),
.X(net579)
);

sky130_fd_sc_hd__mux4_2 c715(
.A0(net577),
.A1(net328),
.A2(net576),
.A3(net474),
.S0(net824),
.S1(net852),
.X(net580)
);

sky130_fd_sc_hd__mux4_1 c716(
.A0(net561),
.A1(net104),
.A2(net528),
.A3(net571),
.S0(net849),
.S1(net851),
.X(net581)
);

sky130_fd_sc_hd__mux4_2 c717(
.A0(net576),
.A1(in46),
.A2(net751),
.A3(net824),
.S0(net842),
.S1(net852),
.X(net582)
);

sky130_fd_sc_hd__mux4_2 c718(
.A0(net554),
.A1(net571),
.A2(net568),
.A3(net842),
.S0(net847),
.S1(net852),
.X(net583)
);

sky130_fd_sc_hd__mux4_1 c719(
.A0(net474),
.A1(net528),
.A2(net846),
.A3(net848),
.S0(net850),
.S1(net854),
.X(net584)
);

sky130_fd_sc_hd__mux4_2 c720(
.A0(net422),
.A1(net372),
.A2(net706),
.A3(net749),
.S0(net849),
.S1(net851),
.X(net585)
);

sky130_fd_sc_hd__mux4_4 c721(
.A0(net547),
.A1(in0),
.A2(net585),
.A3(net751),
.S0(net845),
.S1(net854),
.X(net586)
);

sky130_fd_sc_hd__mux4_4 c722(
.A0(net422),
.A1(net585),
.A2(net122),
.A3(net554),
.S0(net113),
.S1(net841),
.X(net587)
);

sky130_fd_sc_hd__mux4_1 c723(
.A0(net568),
.A1(net586),
.A2(net547),
.A3(net751),
.S0(net842),
.S1(net851),
.X(net588)
);

sky130_fd_sc_hd__mux4_2 c724(
.A0(net474),
.A1(net576),
.A2(net541),
.A3(net699),
.S0(net720),
.S1(net854),
.X(net589)
);

sky130_fd_sc_hd__mux4_2 c725(
.A0(net571),
.A1(net474),
.A2(net720),
.A3(net751),
.S0(net842),
.S1(net854),
.X(net590)
);

sky130_fd_sc_hd__mux4_1 c726(
.A0(net237),
.A1(in13),
.A2(net328),
.A3(net813),
.S0(net841),
.S1(net853),
.X(net591)
);

sky130_fd_sc_hd__mux4_2 c727(
.A0(net541),
.A1(net344),
.A2(net542),
.A3(net104),
.S0(net838),
.S1(net842),
.X(net592)
);

sky130_fd_sc_hd__mux4_1 c728(
.A0(net237),
.A1(net698),
.A2(net753),
.A3(net788),
.S0(net850),
.S1(net856),
.X(net593)
);

sky130_fd_sc_hd__mux4_4 c729(
.A0(net592),
.A1(net386),
.A2(net328),
.A3(net483),
.S0(net753),
.S1(net856),
.X(net594)
);

sky130_fd_sc_hd__mux4_2 c730(
.A0(net592),
.A1(net698),
.A2(net844),
.A3(net852),
.S0(net855),
.S1(net857),
.X(net595)
);

sky130_fd_sc_hd__mux4_4 c731(
.A0(net483),
.A1(net344),
.A2(net386),
.A3(net394),
.S0(net556),
.S1(net698),
.X(net596)
);

sky130_fd_sc_hd__mux4_1 c732(
.A0(net592),
.A1(net542),
.A2(net741),
.A3(net754),
.S0(net844),
.S1(net859),
.X(net597)
);

sky130_fd_sc_hd__mux4_2 c733(
.A0(net597),
.A1(net556),
.A2(net455),
.A3(net18),
.S0(net832),
.S1(net856),
.X(net598)
);

sky130_fd_sc_hd__mux4_4 c734(
.A0(net483),
.A1(in13),
.A2(net595),
.A3(net592),
.S0(net788),
.S1(net841),
.X(net599)
);

sky130_fd_sc_hd__mux4_4 c735(
.A0(net344),
.A1(net592),
.A2(net591),
.A3(in2),
.S0(net715),
.S1(net859),
.X(net600)
);

sky130_fd_sc_hd__mux4_2 c736(
.A0(net455),
.A1(net284),
.A2(net725),
.A3(net741),
.S0(net857),
.S1(net860),
.X(net601)
);

sky130_fd_sc_hd__mux4_1 c737(
.A0(net592),
.A1(net595),
.A2(net601),
.A3(net528),
.S0(net542),
.S1(net697),
.X(net602)
);

sky130_fd_sc_hd__mux4_4 c738(
.A0(net386),
.A1(net591),
.A2(net77),
.A3(net716),
.S0(net736),
.S1(net858),
.X(net603)
);

sky130_fd_sc_hd__mux4_1 c739(
.A0(net541),
.A1(net725),
.A2(net736),
.A3(net842),
.S0(net844),
.S1(net853),
.X(net604)
);

sky130_fd_sc_hd__mux4_1 c740(
.A0(net591),
.A1(net344),
.A2(in31),
.A3(net751),
.S0(net832),
.S1(net858),
.X(net605)
);

sky130_fd_sc_hd__mux4_1 c741(
.A0(net113),
.A1(net483),
.A2(net604),
.A3(net542),
.S0(net751),
.S1(net853),
.X(net606)
);

sky130_fd_sc_hd__mux4_1 c742(
.A0(net215),
.A1(net284),
.A2(net328),
.A3(net715),
.S0(net751),
.S1(net837),
.X(net607)
);

sky130_fd_sc_hd__mux4_2 c743(
.A0(net606),
.A1(net18),
.A2(net454),
.A3(net698),
.S0(net736),
.S1(net751),
.X(net608)
);

sky130_fd_sc_hd__mux4_4 c744(
.A0(net528),
.A1(net595),
.A2(net344),
.A3(net604),
.S0(net725),
.S1(net855),
.X(net609)
);

sky130_fd_sc_hd__mux4_1 c745(
.A0(net394),
.A1(net604),
.A2(net607),
.A3(net344),
.S0(net697),
.S1(net852),
.X(net610)
);

sky130_fd_sc_hd__mux4_1 c746(
.A0(net593),
.A1(net604),
.A2(net386),
.A3(net724),
.S0(net853),
.S1(net855),
.X(net611)
);

sky130_fd_sc_hd__mux4_4 c747(
.A0(net601),
.A1(net606),
.A2(net386),
.A3(net698),
.S0(net699),
.S1(net838),
.X(net612)
);

sky130_fd_sc_hd__mux4_2 c748(
.A0(net601),
.A1(net97),
.A2(net115),
.A3(net215),
.S0(net716),
.S1(net741),
.X(net613)
);

sky130_fd_sc_hd__mux4_2 c749(
.A0(net203),
.A1(net122),
.A2(in2),
.A3(net798),
.S0(net840),
.S1(net850),
.X(net614)
);

sky130_fd_sc_hd__mux4_4 c750(
.A0(net542),
.A1(net122),
.A2(net510),
.A3(net372),
.S0(net798),
.S1(net840),
.X(net615)
);

sky130_fd_sc_hd__mux4_4 c751(
.A0(net18),
.A1(net522),
.A2(net724),
.A3(net747),
.S0(net821),
.S1(net860),
.X(net616)
);

sky130_fd_sc_hd__mux4_1 c752(
.A0(in0),
.A1(net614),
.A2(net522),
.A3(net747),
.S0(net846),
.S1(net860),
.X(net617)
);

sky130_fd_sc_hd__mux4_1 c753(
.A0(net617),
.A1(net18),
.A2(net778),
.A3(net813),
.S0(net817),
.S1(net832),
.X(net618)
);

sky130_fd_sc_hd__mux4_4 c754(
.A0(net522),
.A1(net617),
.A2(net736),
.A3(net752),
.S0(net788),
.S1(net850),
.X(net619)
);

sky130_fd_sc_hd__mux4_4 c755(
.A0(in31),
.A1(net510),
.A2(in0),
.A3(net716),
.S0(net752),
.S1(net844),
.X(net620)
);

sky130_fd_sc_hd__mux4_2 c756(
.A0(net510),
.A1(net542),
.A2(net522),
.A3(net455),
.S0(net724),
.S1(net798),
.X(net621)
);

sky130_fd_sc_hd__mux4_4 c757(
.A0(net607),
.A1(net621),
.A2(net752),
.A3(net798),
.S0(net832),
.S1(net844),
.X(net622)
);

sky130_fd_sc_hd__mux4_2 c758(
.A0(net97),
.A1(net284),
.A2(net706),
.A3(net778),
.S0(net813),
.S1(net846),
.X(net623)
);

sky130_fd_sc_hd__mux4_2 c759(
.A0(net284),
.A1(net616),
.A2(net215),
.A3(net483),
.S0(net741),
.S1(net842),
.X(net624)
);

sky130_fd_sc_hd__mux4_4 c760(
.A0(net372),
.A1(net697),
.A2(net736),
.A3(net747),
.S0(net813),
.S1(net840),
.X(net625)
);

sky130_fd_sc_hd__mux4_1 c761(
.A0(net613),
.A1(net18),
.A2(net620),
.A3(net625),
.S0(net752),
.S1(net840),
.X(net626)
);

sky130_fd_sc_hd__mux4_4 c762(
.A0(net623),
.A1(net510),
.A2(net697),
.A3(net716),
.S0(net778),
.S1(net815),
.X(net627)
);

sky130_fd_sc_hd__mux4_1 c763(
.A0(net626),
.A1(net627),
.A2(net736),
.A3(net741),
.S0(net832),
.S1(net837),
.X(net628)
);

sky130_fd_sc_hd__mux4_4 c764(
.A0(net623),
.A1(net615),
.A2(net625),
.A3(net628),
.S0(net115),
.S1(in41),
.X(net629)
);

sky130_fd_sc_hd__a2111o_1 merge765(
.A1(net83),
.A2(net418),
.B1(net419),
.C1(net88),
.D1(net802),
.X(net630)
);

sky130_fd_sc_hd__mux4_2 merge766(
.A0(net31),
.A1(net44),
.A2(in2),
.A3(in51),
.S0(net48),
.S1(net32),
.X(net631)
);

sky130_fd_sc_hd__mux4_4 merge767(
.A0(net419),
.A1(net425),
.A2(net320),
.A3(net78),
.S0(net424),
.S1(net217),
.X(net632)
);

sky130_fd_sc_hd__o2111ai_2 merge768(
.A1(net29),
.A2(net31),
.B1(net28),
.C1(net16),
.D1(net25),
.Y(net633)
);

sky130_fd_sc_hd__o2111ai_4 merge769(
.A1(net240),
.A2(net209),
.B1(net131),
.C1(net644),
.D1(net657),
.Y(net634)
);

sky130_fd_sc_hd__o2111a_4 merge770(
.A1(net77),
.A2(net208),
.B1(net209),
.C1(net82),
.D1(net214),
.X(net635)
);

sky130_fd_sc_hd__a2111oi_1 merge771(
.A1(net420),
.A2(net419),
.B1(net421),
.C1(net76),
.D1(net424),
.Y(net636)
);

sky130_fd_sc_hd__mux4_1 merge772(
.A0(net211),
.A1(net320),
.A2(net203),
.A3(net74),
.S0(net420),
.S1(net425),
.X(net637)
);

sky130_fd_sc_hd__mux4_1 merge773(
.A0(net231),
.A1(out61),
.A2(net246),
.A3(net243),
.S0(net245),
.S1(net131),
.X(net638)
);

sky130_fd_sc_hd__mux4_1 merge774(
.A0(net425),
.A1(net524),
.A2(net419),
.A3(net533),
.S0(net418),
.S1(net700),
.X(net639)
);

sky130_fd_sc_hd__mux4_2 merge775(
.A0(net418),
.A1(net320),
.A2(net81),
.A3(net531),
.S0(net532),
.S1(net528),
.X(net640)
);

sky130_fd_sc_hd__nor2_2 merge776(
.A(net53),
.B(net59),
.Y(net641)
);

sky130_fd_sc_hd__and2_4 merge777(
.A(net176),
.B(net186),
.X(net642)
);

sky130_fd_sc_hd__dfrbp_1 merge778(
.D(net125),
.RESET_B(net126),
.CLK(clk),
.Q(net644),
.Q_N(net643)
);

sky130_fd_sc_hd__nor2b_4 merge779(
.A(net287),
.B_N(net304),
.Y(net645)
);

sky130_fd_sc_hd__nand2_2 merge780(
.A(net509),
.B(net519),
.Y(net646)
);

sky130_fd_sc_hd__and2b_1 merge781(
.A_N(net152),
.B(net139),
.X(net647)
);

sky130_fd_sc_hd__dfrbp_2 merge782(
.D(net319),
.RESET_B(net323),
.CLK(clk),
.Q(net649),
.Q_N(net648)
);

sky130_fd_sc_hd__dfrtn_1 merge783(
.D(net337),
.RESET_B(net338),
.CLK_N(clk),
.Q(net650)
);

sky130_fd_sc_hd__nor2_1 merge784(
.A(net362),
.B(net361),
.Y(net651)
);

sky130_fd_sc_hd__nor2b_1 merge785(
.A(net444),
.B_N(net456),
.Y(net652)
);

sky130_fd_sc_hd__dfrtp_1 merge786(
.D(net553),
.RESET_B(net559),
.CLK(clk),
.Q(net653)
);

sky130_fd_sc_hd__or2_4 merge787(
.A(net109),
.B(net110),
.X(net654)
);

sky130_fd_sc_hd__nor2b_4 merge788(
.A(net472),
.B_N(net480),
.Y(net655)
);

sky130_fd_sc_hd__and2b_1 merge789(
.A_N(net410),
.B(net411),
.X(net656)
);

sky130_fd_sc_hd__dfrtp_2 merge790(
.D(net227),
.Q(net233),
.CLK(clk)
);

sky130_fd_sc_hd__nand2b_2 merge791(
.A_N(net527),
.B(net536),
.Y(net658)
);

sky130_fd_sc_hd__dfrtp_4 merge792(
.Q(net306),
.RESET_B(net305),
.CLK(clk)
);

sky130_fd_sc_hd__nand2_2 merge793(
.A(net437),
.B(net630),
.Y(net659)
);

sky130_fd_sc_hd__and2b_1 merge794(
.A_N(net382),
.B(net398),
.X(net660)
);

sky130_fd_sc_hd__dfsbp_1 merge795(
.D(net283),
.SET_B(net271),
.CLK(clk),
.Q(net662),
.Q_N(net661)
);

sky130_fd_sc_hd__nor2_4 merge796(
.A(net629),
.B(net619),
.Y(net663)
);

sky130_fd_sc_hd__and2_2 merge797(
.A(net491),
.B(net494),
.X(net664)
);

sky130_fd_sc_hd__dfsbp_2 merge798(
.D(net47),
.SET_B(net633),
.CLK(clk),
.Q(net666),
.Q_N(net665)
);

sky130_fd_sc_hd__dfstp_1 merge799(
.D(net163),
.SET_B(net164),
.CLK(clk),
.Q(out47)
);

sky130_fd_sc_hd__nor2b_4 merge800(
.A(net594),
.B_N(net605),
.Y(net667)
);

sky130_fd_sc_hd__dfstp_2 merge801(
.D(net218),
.SET_B(net210),
.CLK(clk),
.Q(net668)
);

sky130_fd_sc_hd__nor2b_2 merge802(
.A(net572),
.B_N(net578),
.Y(net669)
);

sky130_fd_sc_hd__nand2b_4 merge803(
.A_N(net252),
.B(net256),
.Y(net670)
);

sky130_fd_sc_hd__and2b_1 merge804(
.A_N(net460),
.B(net457),
.X(net671)
);

sky130_fd_sc_hd__dfstp_4 merge805(
.D(net374),
.SET_B(net638),
.CLK(clk),
.Q(net672)
);

sky130_fd_sc_hd__dlrbn_1 merge806(
.D(net216),
.RESET_B(net236),
.GATE_N(clk),
.Q(net674),
.Q_N(net673)
);

sky130_fd_sc_hd__dlrbn_2 merge807(
.D(net354),
.RESET_B(net635),
.GATE_N(clk),
.Q(net676),
.Q_N(net675)
);

sky130_fd_sc_hd__or2_4 merge808(
.A(net413),
.B(net417),
.X(net677)
);

sky130_fd_sc_hd__or2b_1 merge809(
.A(net482),
.B_N(net520),
.X(net678)
);

sky130_fd_sc_hd__and2b_4 merge810(
.A_N(net142),
.B(net143),
.X(net679)
);

sky130_fd_sc_hd__dlrbp_1 merge811(
.D(net151),
.RESET_B(net154),
.GATE(clk),
.Q(net681),
.Q_N(net680)
);

sky130_fd_sc_hd__dlrbp_2 merge812(
.D(net664),
.RESET_B(net502),
.GATE(clk),
.Q(net683),
.Q_N(net682)
);

sky130_fd_sc_hd__dlrtn_1 merge813(
.D(net352),
.RESET_B(net655),
.GATE_N(clk),
.Q(net684)
);

sky130_fd_sc_hd__dlrtn_2 merge814(
.D(net652),
.RESET_B(net449),
.GATE_N(clk),
.Q(net685)
);

sky130_fd_sc_hd__or2b_4 merge815(
.A(net584),
.B_N(net622),
.X(net686)
);

sky130_fd_sc_hd__nor2_2 merge816(
.A(net663),
.B(net646),
.Y(net687)
);

sky130_fd_sc_hd__nand2_4 merge817(
.A(net588),
.B(net611),
.Y(net688)
);

sky130_fd_sc_hd__nand2b_4 merge818(
.A_N(net416),
.B(net290),
.Y(net689)
);

sky130_fd_sc_hd__nand2_2 merge819(
.A(net642),
.B(net63),
.Y(net690)
);

sky130_fd_sc_hd__and2b_1 merge820(
.A_N(net387),
.B(net293),
.X(net691)
);

sky130_fd_sc_hd__nand2_2 merge821(
.A(net609),
.B(net598),
.Y(net692)
);

sky130_fd_sc_hd__nand2_4 merge822(
.A(net193),
.B(net631),
.Y(net693)
);

sky130_fd_sc_hd__and2_4 merge823(
.A(net589),
.B(net570),
.X(net694)
);

sky130_fd_sc_hd__nor2b_2 merge824(
.A(net167),
.B_N(net150),
.Y(net695)
);

sky130_fd_sc_hd__dlrtn_4 merge825(
.D(net632),
.RESET_B(net658),
.GATE_N(clk),
.Q(net696)
);

sky130_fd_sc_hd__dlrtp_1 merge826(
.D(net600),
.RESET_B(net624),
.GATE(clk),
.Q(net697)
);

sky130_fd_sc_hd__dlrtp_2 merge827(
.D(net654),
.RESET_B(net111),
.GATE(clk),
.Q(net698)
);

sky130_fd_sc_hd__dlrtp_4 merge828(
.D(net370),
.RESET_B(net677),
.GATE(clk),
.Q(out40)
);

sky130_fd_sc_hd__edfxbp_1 merge829(
.D(net538),
.DE(net688),
.CLK(clk),
.Q(net700),
.Q_N(net699)
);

sky130_fd_sc_hd__or2_2 merge830(
.A(net660),
.B(net656),
.X(net701)
);

sky130_fd_sc_hd__edfxtp_1 merge831(
.D(net41),
.DE(net195),
.CLK(clk),
.Q(net702)
);

sky130_fd_sc_hd__nand2_1 merge832(
.A(net258),
.B(net299),
.Y(net703)
);

sky130_fd_sc_hd__or2b_4 merge833(
.A(net634),
.B_N(net388),
.X(net704)
);

sky130_fd_sc_hd__sdlclkp_1 merge834(
.GATE(net406),
.SCE(net402),
.CLK(clk),
.GCLK(out30)
);

sky130_fd_sc_hd__sdlclkp_2 merge835(
.GATE(net645),
.SCE(net647),
.CLK(clk),
.GCLK(net705)
);

sky130_fd_sc_hd__sdlclkp_4 merge836(
.GATE(net636),
.SCE(net686),
.CLK(clk),
.GCLK(net706)
);

sky130_fd_sc_hd__and2_2 merge837(
.A(net670),
.B(net260),
.X(net707)
);

sky130_fd_sc_hd__dfrbp_1 merge838(
.D(net132),
.Q(net709),
.CLK(clk),
.Q_N(net708)
);

sky130_fd_sc_hd__or2_2 merge839(
.A(net379),
.B(net385),
.X(net710)
);

sky130_fd_sc_hd__or2_4 merge840(
.A(net651),
.B(net669),
.X(net711)
);

sky130_fd_sc_hd__nor2_1 merge841(
.A(net383),
.B(net384),
.Y(net712)
);

sky130_fd_sc_hd__dfrbp_2 merge842(
.D(net313),
.RESET_B(net367),
.CLK(clk),
.Q(net714),
.Q_N(net713)
);

sky130_fd_sc_hd__dfrtn_1 merge843(
.D(net667),
.RESET_B(net468),
.CLK_N(clk),
.Q(net715)
);

sky130_fd_sc_hd__dfrtp_1 merge844(
.D(net687),
.RESET_B(net596),
.CLK(clk),
.Q(net716)
);

sky130_fd_sc_hd__dfrtp_2 merge845(
.D(net678),
.RESET_B(net476),
.CLK(clk),
.Q(net717)
);

sky130_fd_sc_hd__nor2_2 merge846(
.A(net637),
.B(net477),
.Y(net718)
);

sky130_fd_sc_hd__dfrtp_4 merge847(
.D(net640),
.RESET_B(net639),
.CLK(clk),
.Q(net719)
);

sky130_fd_sc_hd__dfsbp_1 merge848(
.D(net488),
.SET_B(net694),
.CLK(clk),
.Q(net721),
.Q_N(net720)
);

sky130_fd_sc_hd__dfsbp_2 merge849(
.D(net432),
.SET_B(net518),
.CLK(clk),
.Q(net723),
.Q_N(net722)
);

sky130_fd_sc_hd__dfstp_1 merge850(
.D(net692),
.SET_B(net479),
.CLK(clk),
.Q(net724)
);

sky130_fd_sc_hd__dfstp_2 merge851(
.D(net689),
.SET_B(net599),
.CLK(clk),
.Q(net725)
);

sky130_fd_sc_hd__dfstp_4 merge852(
.D(net427),
.SET_B(net671),
.CLK(clk),
.Q(net726)
);

sky130_fd_sc_hd__dlrbn_1 merge853(
.D(net537),
.RESET_B(net279),
.GATE_N(clk),
.Q(net728),
.Q_N(net727)
);

sky130_fd_sc_hd__dlrbn_2 merge854(
.D(net436),
.RESET_B(net565),
.GATE_N(clk),
.Q(net730),
.Q_N(net729)
);

sky130_fd_sc_hd__dlrbp_1 merge855(
.D(net178),
.RESET_B(net489),
.GATE(clk),
.Q(net732),
.Q_N(net731)
);

sky130_fd_sc_hd__dlrbp_2 merge856(
.D(net703),
.RESET_B(net278),
.GATE(clk),
.Q(net734),
.Q_N(net733)
);

sky130_fd_sc_hd__dlrtn_1 merge857(
.D(net414),
.RESET_B(net405),
.GATE_N(clk),
.Q(net735)
);

sky130_fd_sc_hd__dlrtn_2 merge858(
.D(net612),
.RESET_B(net602),
.GATE_N(clk),
.Q(net736)
);

sky130_fd_sc_hd__dlrtn_4 merge859(
.D(net695),
.RESET_B(net294),
.GATE_N(clk),
.Q(out48)
);

sky130_fd_sc_hd__dlrtp_1 merge860(
.D(net189),
.RESET_B(net641),
.GATE(clk),
.Q(out36)
);

sky130_fd_sc_hd__dlrtp_2 merge861(
.D(net659),
.RESET_B(net718),
.GATE(clk),
.Q(net737)
);

sky130_fd_sc_hd__dlrtp_4 merge862(
.D(net704),
.RESET_B(net710),
.GATE(clk),
.Q(net738)
);

sky130_fd_sc_hd__edfxbp_1 merge863(
.Q_N(net266),
.DE(net263),
.CLK(clk),
.Q(net740)
);

sky130_fd_sc_hd__edfxtp_1 merge864(
.D(net546),
.DE(net610),
.CLK(clk),
.Q(net741)
);

sky130_fd_sc_hd__sdlclkp_1 merge865(
.GATE(net539),
.SCE(net550),
.CLK(clk),
.GCLK(net742)
);

sky130_fd_sc_hd__sdlclkp_2 merge866(
.GATE(net148),
.SCE(net693),
.CLK(clk),
.GCLK(net743)
);

sky130_fd_sc_hd__sdlclkp_4 merge867(
.GATE(net679),
.SCE(net690),
.CLK(clk),
.GCLK(net744)
);

sky130_fd_sc_hd__dfrbp_1 merge868(
.D(net269),
.RESET_B(net291),
.CLK(clk),
.Q(net746),
.Q_N(net745)
);

sky130_fd_sc_hd__dfrbp_2 merge869(
.D(net549),
.RESET_B(net608),
.CLK(clk),
.Q(net748),
.Q_N(net747)
);

sky130_fd_sc_hd__dfrtn_1 merge870(
.D(net711),
.RESET_B(net180),
.CLK_N(clk),
.Q(net749)
);

sky130_fd_sc_hd__dfrtp_1 merge871(
.D(net114),
.RESET_B(net707),
.CLK(clk),
.Q(net750)
);

sky130_fd_sc_hd__dfrtp_2 merge872(
.D(net691),
.RESET_B(net701),
.CLK(clk),
.Q(out49)
);

sky130_fd_sc_hd__dfrtp_4 merge873(
.D(net603),
.RESET_B(net581),
.CLK(clk),
.Q(net751)
);

sky130_fd_sc_hd__dfsbp_1 merge874(
.D(net712),
.SET_B(net618),
.CLK(clk),
.Q(out42),
.Q_N(net752)
);

sky130_fd_sc_hd__dfsbp_2 merge875(
.D(net564),
.SET_B(net540),
.CLK(clk),
.Q(net754),
.Q_N(net753)
);

sky130_fd_sc_hd__dfxbp_1 s876(
.D(net43),
.CLK(clk),
.Q(net756),
.Q_N(net755)
);

sky130_fd_sc_hd__dfxbp_2 s877(
.D(net108),
.CLK(clk),
.Q(net758),
.Q_N(net757)
);

sky130_fd_sc_hd__dfxtp_1 s878(
.D(net120),
.CLK(clk),
.Q(out5)
);

sky130_fd_sc_hd__dfxtp_2 s879(
.D(net144),
.CLK(clk),
.Q(net759)
);

sky130_fd_sc_hd__dfxtp_4 s880(
.D(net155),
.CLK(clk),
.Q(out52)
);

sky130_fd_sc_hd__dlclkp_1 s881(
.GATE(net156),
.CLK(clk),
.GCLK(net760)
);

sky130_fd_sc_hd__dlclkp_2 s882(
.GATE(net157),
.CLK(clk),
.GCLK(net761)
);

sky130_fd_sc_hd__dlclkp_4 s883(
.GATE(net158),
.CLK(clk),
.GCLK(net762)
);

sky130_fd_sc_hd__dlxbn_1 s884(
.D(net159),
.GATE_N(clk),
.Q(net764),
.Q_N(net763)
);

sky130_fd_sc_hd__dlxbn_2 s885(
.D(net160),
.GATE_N(clk),
.Q(out15),
.Q_N(net765)
);

sky130_fd_sc_hd__dlxbp_1 s886(
.D(net161),
.GATE(clk),
.Q(net767),
.Q_N(net766)
);

sky130_fd_sc_hd__dlxtn_1 s887(
.D(net162),
.GATE_N(clk),
.Q(net768)
);

sky130_fd_sc_hd__dlxtn_2 s888(
.D(net165),
.GATE_N(clk),
.Q(net769)
);

sky130_fd_sc_hd__dlxtn_4 s889(
.D(net166),
.GATE_N(clk),
.Q(net770)
);

sky130_fd_sc_hd__dlxtp_1 s890(
.D(net170),
.GATE(clk),
.Q(net771)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s891(
.D(net173),
.SLEEP_B(clk),
.Q(net772)
);

sky130_fd_sc_hd__dfxbp_1 s892(
.D(net183),
.CLK(clk),
.Q(out43),
.Q_N(net773)
);

sky130_fd_sc_hd__dfxbp_2 s893(
.D(net187),
.CLK(clk),
.Q(net775),
.Q_N(net774)
);

sky130_fd_sc_hd__dfxtp_1 s894(
.D(net190),
.CLK(clk),
.Q(net776)
);

sky130_fd_sc_hd__dfxtp_2 s895(
.D(net219),
.CLK(clk),
.Q(net777)
);

sky130_fd_sc_hd__dfxtp_4 s896(
.D(net226),
.CLK(clk),
.Q(out1)
);

sky130_fd_sc_hd__dlclkp_1 s897(
.GATE(net235),
.CLK(clk),
.GCLK(net778)
);

sky130_fd_sc_hd__dlclkp_2 s898(
.GATE(net239),
.CLK(clk),
.GCLK(net779)
);

sky130_fd_sc_hd__dlclkp_4 s899(
.GATE(net244),
.CLK(clk),
.GCLK(net780)
);

sky130_fd_sc_hd__dlxbn_1 s900(
.D(net248),
.GATE_N(clk),
.Q(net782),
.Q_N(net781)
);

sky130_fd_sc_hd__dlxbn_2 s901(
.D(net259),
.GATE_N(clk),
.Q(out7),
.Q_N(net783)
);

sky130_fd_sc_hd__dlxbp_1 s902(
.D(net262),
.GATE(clk),
.Q(net785),
.Q_N(net784)
);

sky130_fd_sc_hd__dlxtn_1 s903(
.D(net264),
.GATE_N(clk),
.Q(net786)
);

sky130_fd_sc_hd__dlxtn_2 s904(
.D(net265),
.GATE_N(clk),
.Q(net787)
);

sky130_fd_sc_hd__dlxtn_4 s905(
.D(net267),
.GATE_N(clk),
.Q(net788)
);

sky130_fd_sc_hd__dlxtp_1 s906(
.D(net268),
.GATE(clk),
.Q(net789)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s907(
.D(net270),
.SLEEP_B(clk),
.Q(net790)
);

sky130_fd_sc_hd__dfxbp_1 s908(
.D(net274),
.CLK(clk),
.Q(out56),
.Q_N(net791)
);

sky130_fd_sc_hd__dfxbp_2 s909(
.D(net276),
.CLK(clk),
.Q(net793),
.Q_N(net792)
);

sky130_fd_sc_hd__dfxtp_1 s910(
.D(net277),
.CLK(clk),
.Q(net794)
);

sky130_fd_sc_hd__dfxtp_2 s911(
.D(net280),
.CLK(clk),
.Q(net795)
);

sky130_fd_sc_hd__dfxtp_4 s912(
.D(net286),
.CLK(clk),
.Q(net796)
);

sky130_fd_sc_hd__dlclkp_1 s913(
.GATE(net298),
.CLK(clk),
.GCLK(net797)
);

sky130_fd_sc_hd__dlclkp_2 s914(
.GATE(net301),
.CLK(clk),
.GCLK(net798)
);

sky130_fd_sc_hd__dlclkp_4 s915(
.GATE(net325),
.CLK(clk),
.GCLK(net799)
);

sky130_fd_sc_hd__dlxbn_1 s916(
.D(net326),
.GATE_N(clk),
.Q(net801),
.Q_N(net800)
);

sky130_fd_sc_hd__dlxbn_2 s917(
.D(net327),
.GATE_N(clk),
.Q(net803),
.Q_N(net802)
);

sky130_fd_sc_hd__dlxbp_1 s918(
.D(net336),
.GATE(clk),
.Q(net805),
.Q_N(net804)
);

sky130_fd_sc_hd__dlxtn_1 s919(
.D(net349),
.GATE_N(clk),
.Q(net806)
);

sky130_fd_sc_hd__dlxtn_2 s920(
.D(net350),
.GATE_N(clk),
.Q(out24)
);

sky130_fd_sc_hd__dlxtn_4 s921(
.D(net353),
.GATE_N(clk),
.Q(net807)
);

sky130_fd_sc_hd__dlxtp_1 s922(
.D(net355),
.GATE(clk),
.Q(net808)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s923(
.D(net380),
.SLEEP_B(clk),
.Q(out39)
);

sky130_fd_sc_hd__dfxbp_1 s924(
.D(net381),
.CLK(clk),
.Q(net810),
.Q_N(net809)
);

sky130_fd_sc_hd__dfxbp_2 s925(
.D(net389),
.CLK(clk),
.Q(net812),
.Q_N(net811)
);

sky130_fd_sc_hd__dfxtp_1 s926(
.D(net392),
.CLK(clk),
.Q(out9)
);

sky130_fd_sc_hd__dfxtp_2 s927(
.D(net395),
.CLK(clk),
.Q(net813)
);

sky130_fd_sc_hd__dfxtp_4 s928(
.D(net399),
.CLK(clk),
.Q(net814)
);

sky130_fd_sc_hd__dlclkp_1 s929(
.GATE(net404),
.CLK(clk),
.GCLK(out13)
);

sky130_fd_sc_hd__dlclkp_2 s930(
.GATE(net407),
.CLK(clk),
.GCLK(net815)
);

sky130_fd_sc_hd__dlclkp_4 s931(
.GATE(net408),
.CLK(clk),
.GCLK(out10)
);

sky130_fd_sc_hd__dlxbn_1 s932(
.D(net409),
.GATE_N(clk),
.Q(net817),
.Q_N(net816)
);

sky130_fd_sc_hd__dlxbn_2 s933(
.D(net412),
.GATE_N(clk),
.Q(net819),
.Q_N(net818)
);

sky130_fd_sc_hd__dlxbp_1 s934(
.D(net415),
.GATE(clk),
.Q(net821),
.Q_N(net820)
);

sky130_fd_sc_hd__dlxtn_1 s935(
.D(net434),
.GATE_N(clk),
.Q(net822)
);

sky130_fd_sc_hd__dlxtn_2 s936(
.D(net435),
.GATE_N(clk),
.Q(net823)
);

sky130_fd_sc_hd__dlxtn_4 s937(
.D(net438),
.GATE_N(clk),
.Q(net824)
);

sky130_fd_sc_hd__dlxtp_1 s938(
.D(net458),
.GATE(clk),
.Q(net825)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s939(
.D(net459),
.SLEEP_B(clk),
.Q(out21)
);

sky130_fd_sc_hd__dfxbp_1 s940(
.D(net463),
.CLK(clk),
.Q(net827),
.Q_N(net826)
);

sky130_fd_sc_hd__dfxbp_2 s941(
.D(net466),
.CLK(clk),
.Q(net829),
.Q_N(net828)
);

sky130_fd_sc_hd__dfxtp_1 s942(
.D(net470),
.CLK(clk),
.Q(net830)
);

sky130_fd_sc_hd__dfxtp_2 s943(
.D(net473),
.CLK(clk),
.Q(net831)
);

sky130_fd_sc_hd__dfxtp_4 s944(
.D(net478),
.CLK(clk),
.Q(net832)
);

sky130_fd_sc_hd__dlclkp_1 s945(
.GATE(net495),
.CLK(clk),
.GCLK(net833)
);

sky130_fd_sc_hd__dlclkp_2 s946(
.GATE(net496),
.CLK(clk),
.GCLK(net834)
);

sky130_fd_sc_hd__dlclkp_4 s947(
.GATE(net497),
.CLK(clk),
.GCLK(net835)
);

sky130_fd_sc_hd__dlxbn_1 s948(
.D(net501),
.GATE_N(clk),
.Q(out19),
.Q_N(net836)
);

sky130_fd_sc_hd__dlxbn_2 s949(
.D(net503),
.GATE_N(clk),
.Q(net838),
.Q_N(net837)
);

sky130_fd_sc_hd__dlxbp_1 s950(
.D(net504),
.GATE(clk),
.Q(out3),
.Q_N(net839)
);

sky130_fd_sc_hd__dlxtn_1 s951(
.D(net523),
.GATE_N(clk),
.Q(net840)
);

sky130_fd_sc_hd__dlxtn_2 s952(
.D(net534),
.GATE_N(clk),
.Q(net841)
);

sky130_fd_sc_hd__dlxtn_4 s953(
.D(net545),
.GATE_N(clk),
.Q(net842)
);

sky130_fd_sc_hd__dlxtp_1 s954(
.D(net563),
.GATE(clk),
.Q(net843)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s955(
.D(net566),
.SLEEP_B(clk),
.Q(net844)
);

sky130_fd_sc_hd__dfxbp_1 s956(
.D(net567),
.CLK(clk),
.Q(net846),
.Q_N(net845)
);

sky130_fd_sc_hd__dfxbp_2 s957(
.D(net569),
.CLK(clk),
.Q(net848),
.Q_N(net847)
);

sky130_fd_sc_hd__dfxtp_1 s958(
.D(net573),
.CLK(clk),
.Q(net849)
);

sky130_fd_sc_hd__dfxtp_2 s959(
.D(net574),
.CLK(clk),
.Q(net850)
);

sky130_fd_sc_hd__dfxtp_4 s960(
.D(net575),
.CLK(clk),
.Q(net851)
);

sky130_fd_sc_hd__dlclkp_1 s961(
.GATE(net579),
.CLK(clk),
.GCLK(net852)
);

sky130_fd_sc_hd__dlclkp_2 s962(
.GATE(net580),
.CLK(clk),
.GCLK(net853)
);

sky130_fd_sc_hd__dlclkp_4 s963(
.GATE(net582),
.CLK(clk),
.GCLK(net854)
);

sky130_fd_sc_hd__dlxbn_1 s964(
.D(net583),
.GATE_N(clk),
.Q(net856),
.Q_N(net855)
);

sky130_fd_sc_hd__dlxbn_2 s965(
.D(net587),
.GATE_N(clk),
.Q(net858),
.Q_N(net857)
);

sky130_fd_sc_hd__dlxbp_1 s966(
.D(net590),
.GATE(clk),
.Q(net860),
.Q_N(net859)
);


endmodule
