module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire clknet_0_clk;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net984;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net635;
 wire net692;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net985;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net802;
 wire clknet_1_0__leaf_net802;
 wire clknet_1_1__leaf_net802;
 wire clknet_0_net370;
 wire clknet_1_0__leaf_net370;
 wire clknet_1_1__leaf_net370;
 wire clknet_0_net381;
 wire clknet_1_0__leaf_net381;
 wire clknet_1_1__leaf_net381;
 wire clknet_0_net704;
 wire clknet_1_0__leaf_net704;
 wire clknet_1_1__leaf_net704;
 wire clknet_0_net409;
 wire clknet_1_0__leaf_net409;
 wire clknet_1_1__leaf_net409;
 wire clknet_0_net705;
 wire clknet_1_0__leaf_net705;
 wire clknet_1_1__leaf_net705;
 wire clknet_0_net780;
 wire clknet_1_0__leaf_net780;
 wire clknet_1_1__leaf_net780;
 wire clknet_0_net625;
 wire clknet_1_0__leaf_net625;
 wire clknet_1_1__leaf_net625;
 wire clknet_0_net626;
 wire clknet_1_0__leaf_net626;
 wire clknet_1_1__leaf_net626;
 wire clknet_0_net703;
 wire clknet_1_0__leaf_net703;
 wire clknet_1_1__leaf_net703;
 wire clknet_0_net628;
 wire clknet_1_0__leaf_net628;
 wire clknet_1_1__leaf_net628;
 wire clknet_0_net616;
 wire clknet_1_0__leaf_net616;
 wire clknet_1_1__leaf_net616;
 wire clknet_0_net880;
 wire clknet_1_0__leaf_net880;
 wire clknet_1_1__leaf_net880;
 wire clknet_0_net386;
 wire clknet_1_0__leaf_net386;
 wire clknet_1_1__leaf_net386;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net779;
 wire clknet_1_0__leaf_net779;
 wire clknet_1_1__leaf_net779;
 wire clknet_0_net876;
 wire clknet_1_0__leaf_net876;
 wire clknet_1_1__leaf_net876;
 wire clknet_0_net490;
 wire clknet_1_0__leaf_net490;
 wire clknet_1_1__leaf_net490;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net403;
 wire clknet_1_0__leaf_net403;
 wire clknet_1_1__leaf_net403;
 wire clknet_0_net385;
 wire clknet_1_0__leaf_net385;
 wire clknet_1_1__leaf_net385;
 wire clknet_0_net901;
 wire clknet_1_0__leaf_net901;
 wire clknet_1_1__leaf_net901;
 wire clknet_0_net893;
 wire clknet_1_0__leaf_net893;
 wire clknet_1_1__leaf_net893;
 wire clknet_0_net906;
 wire clknet_1_0__leaf_net906;
 wire clknet_1_1__leaf_net906;
 wire clknet_0_net911;
 wire clknet_1_0__leaf_net911;
 wire clknet_1_1__leaf_net911;
 wire clknet_0_net482;
 wire clknet_1_0__leaf_net482;
 wire clknet_1_1__leaf_net482;
 wire clknet_0_net397;
 wire clknet_1_0__leaf_net397;
 wire clknet_1_1__leaf_net397;
 wire clknet_0_net618;
 wire clknet_1_0__leaf_net618;
 wire clknet_1_1__leaf_net618;
 wire clknet_0_net382;
 wire clknet_1_0__leaf_net382;
 wire clknet_1_1__leaf_net382;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net801;
 wire clknet_1_0__leaf_net801;
 wire clknet_1_1__leaf_net801;
 wire clknet_0_net467;
 wire clknet_1_0__leaf_net467;
 wire clknet_1_1__leaf_net467;
 wire clknet_0_net569;
 wire clknet_1_0__leaf_net569;
 wire clknet_1_1__leaf_net569;
 wire clknet_0_net581;
 wire clknet_1_0__leaf_net581;
 wire clknet_1_1__leaf_net581;
 wire clknet_0_net583;
 wire clknet_1_0__leaf_net583;
 wire clknet_1_1__leaf_net583;
 wire clknet_0_net800;
 wire clknet_1_0__leaf_net800;
 wire clknet_1_1__leaf_net800;
 wire clknet_0_net471;
 wire clknet_1_0__leaf_net471;
 wire clknet_1_1__leaf_net471;
 wire clknet_0_net474;
 wire clknet_1_0__leaf_net474;
 wire clknet_1_1__leaf_net474;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net249;
 wire clknet_1_0__leaf_net249;
 wire clknet_1_1__leaf_net249;
 wire clknet_0_net781;
 wire clknet_1_0__leaf_net781;
 wire clknet_1_1__leaf_net781;
 wire clknet_0_net557;
 wire clknet_1_0__leaf_net557;
 wire clknet_1_1__leaf_net557;
 wire clknet_0_net558;
 wire clknet_1_0__leaf_net558;
 wire clknet_1_1__leaf_net558;
 wire clknet_0_net575;
 wire clknet_1_0__leaf_net575;
 wire clknet_1_1__leaf_net575;
 wire clknet_0_net568;
 wire clknet_1_0__leaf_net568;
 wire clknet_1_1__leaf_net568;
 wire clknet_0_net560;
 wire clknet_1_0__leaf_net560;
 wire clknet_1_1__leaf_net560;
 wire clknet_0_net761;
 wire clknet_1_0__leaf_net761;
 wire clknet_1_1__leaf_net761;
 wire clknet_0_net760;
 wire clknet_1_0__leaf_net760;
 wire clknet_1_1__leaf_net760;
 wire clknet_0_net759;
 wire clknet_1_0__leaf_net759;
 wire clknet_1_1__leaf_net759;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net453;
 wire clknet_1_0__leaf_net453;
 wire clknet_1_1__leaf_net453;
 wire clknet_0_net551;
 wire clknet_1_0__leaf_net551;
 wire clknet_1_1__leaf_net551;
 wire clknet_0_net450;
 wire clknet_1_0__leaf_net450;
 wire clknet_1_1__leaf_net450;
 wire clknet_0_net552;
 wire clknet_1_0__leaf_net552;
 wire clknet_1_1__leaf_net552;
 wire clknet_0_net744;
 wire clknet_1_0__leaf_net744;
 wire clknet_1_1__leaf_net744;
 wire clknet_0_net371;
 wire clknet_1_0__leaf_net371;
 wire clknet_1_1__leaf_net371;
 wire clknet_0_net322;
 wire clknet_1_0__leaf_net322;
 wire clknet_1_1__leaf_net322;
 wire clknet_0_net743;
 wire clknet_1_0__leaf_net743;
 wire clknet_1_1__leaf_net743;
 wire clknet_0_net317;
 wire clknet_1_0__leaf_net317;
 wire clknet_1_1__leaf_net317;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net908;
 wire clknet_1_0__leaf_net908;
 wire clknet_1_1__leaf_net908;
 wire clknet_0_net727;
 wire clknet_1_0__leaf_net727;
 wire clknet_1_1__leaf_net727;
 wire clknet_0_net151;
 wire clknet_1_0__leaf_net151;
 wire clknet_1_1__leaf_net151;
 wire clknet_0_net153;
 wire clknet_1_0__leaf_net153;
 wire clknet_1_1__leaf_net153;
 wire clknet_0_net152;
 wire clknet_1_0__leaf_net152;
 wire clknet_1_1__leaf_net152;
 wire clknet_0_net261;
 wire clknet_1_0__leaf_net261;
 wire clknet_1_1__leaf_net261;
 wire clknet_0_net147;
 wire clknet_1_0__leaf_net147;
 wire clknet_1_1__leaf_net147;
 wire clknet_0_net726;
 wire clknet_1_0__leaf_net726;
 wire clknet_1_1__leaf_net726;
 wire clknet_0_net465;
 wire clknet_1_0__leaf_net465;
 wire clknet_1_1__leaf_net465;
 wire clknet_0_net459;
 wire clknet_1_0__leaf_net459;
 wire clknet_1_1__leaf_net459;
 wire clknet_0_net350;
 wire clknet_1_0__leaf_net350;
 wire clknet_1_1__leaf_net350;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net245;
 wire clknet_1_0__leaf_net245;
 wire clknet_1_1__leaf_net245;
 wire clknet_0_net252;
 wire clknet_1_0__leaf_net252;
 wire clknet_1_1__leaf_net252;
 wire clknet_0_net247;
 wire clknet_1_0__leaf_net247;
 wire clknet_1_1__leaf_net247;
 wire clknet_0_net130;
 wire clknet_1_0__leaf_net130;
 wire clknet_1_1__leaf_net130;
 wire clknet_0_net725;
 wire clknet_1_0__leaf_net725;
 wire clknet_1_1__leaf_net725;
 wire net363;
 wire net587;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;

 sky130_fd_sc_hd__or2_2 c100 (.A(net36),
    .B(net33),
    .X(net37));
 sky130_fd_sc_hd__nor2_2 c101 (.A(net11),
    .B(net35),
    .Y(net38));
 sky130_fd_sc_hd__nand4_2 c102 (.A(net34),
    .B(net833),
    .C(net38),
    .D(net27),
    .Y(net39));
 sky130_fd_sc_hd__nand4_1 c103 (.A(net29),
    .B(net31),
    .C(net38),
    .D(net27),
    .Y(net40));
 sky130_fd_sc_hd__nand2b_2 c104 (.A_N(net35),
    .B(net38),
    .Y(net41));
 sky130_fd_sc_hd__nor4b_4 c105 (.A(net41),
    .B(net31),
    .C(net38),
    .D_N(net34),
    .Y(net42));
 sky130_fd_sc_hd__mux4_2 c106 (.A0(net32),
    .A1(net36),
    .A2(net5),
    .A3(net26),
    .S0(net861),
    .S1(net41),
    .X(net43));
 sky130_fd_sc_hd__a2111oi_1 c107 (.A1(net40),
    .A2(net43),
    .B1(net41),
    .C1(net891),
    .D1(net42),
    .Y(net44));
 sky130_fd_sc_hd__a2111o_1 c108 (.A1(net37),
    .A2(net1024),
    .B1(net38),
    .C1(net41),
    .D1(net10),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net846),
    .A1(net22),
    .A2(net32),
    .A3(net45),
    .S0(net9),
    .S1(net976),
    .X(net46));
 sky130_fd_sc_hd__nand2_2 c110 (.A(net866),
    .B(net10),
    .Y(net47));
 sky130_fd_sc_hd__nor2b_1 c111 (.A(net946),
    .B_N(net46),
    .Y(net48));
 sky130_fd_sc_hd__and2b_2 c112 (.A_N(net10),
    .B(net30),
    .X(net49));
 sky130_fd_sc_hd__and2b_2 c113 (.A_N(net49),
    .B(net866),
    .X(net50));
 sky130_fd_sc_hd__and2b_1 c114 (.A_N(net47),
    .B(net947),
    .X(net51));
 sky130_fd_sc_hd__and2_2 c115 (.A(net818),
    .B(net27),
    .X(net52));
 sky130_fd_sc_hd__and2b_1 c116 (.A_N(net835),
    .B(net28),
    .X(net53));
 sky130_fd_sc_hd__or2b_1 c117 (.A(net28),
    .B_N(net947),
    .X(net913));
 sky130_fd_sc_hd__and2_2 c118 (.A(net45),
    .B(net10),
    .X(net54));
 sky130_fd_sc_hd__o2111ai_4 c119 (.A1(net48),
    .A2(net842),
    .B1(net947),
    .C1(net47),
    .D1(net49),
    .Y(net55));
 sky130_fd_sc_hd__sdfbbn_1 c120 (.CLK_N(clknet_4_10_0_clk),
    .D(net53),
    .RESET_B(net49),
    .SCD(net55),
    .SCE(net835),
    .SET_B(net27),
    .Q(net57),
    .Q_N(net56));
 sky130_fd_sc_hd__sdfbbn_1 c121 (.CLK_N(clknet_4_10_0_clk),
    .D(net54),
    .RESET_B(net49),
    .SCD(net947),
    .SCE(net838),
    .SET_B(net55),
    .Q(net59),
    .Q_N(net58));
 sky130_fd_sc_hd__nand3b_1 c122 (.A_N(net51),
    .B(net48),
    .C(net58),
    .Y(net60));
 sky130_fd_sc_hd__clkbuf_2 c123 (.A(net902),
    .X(net61));
 sky130_fd_sc_hd__and4b_2 c124 (.A_N(net54),
    .B(net51),
    .C(net46),
    .D(net52),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net16),
    .A1(net59),
    .A2(net62),
    .A3(net60),
    .S0(net49),
    .S1(net47),
    .X(net63));
 sky130_fd_sc_hd__a2111oi_2 c126 (.A1(net59),
    .A2(net52),
    .B1(net61),
    .C1(net62),
    .D1(net719),
    .Y(net64));
 sky130_fd_sc_hd__and2_1 c127 (.A(net47),
    .B(net49),
    .X(net65));
 sky130_fd_sc_hd__a2111oi_1 c128 (.A1(net62),
    .A2(net65),
    .B1(net54),
    .C1(net49),
    .D1(net720),
    .Y(net914));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net30),
    .A1(net847),
    .A2(net53),
    .A3(net861),
    .S0(net64),
    .S1(net719),
    .X(net66));
 sky130_fd_sc_hd__a2111oi_1 c130 (.A1(net64),
    .A2(net1020),
    .B1(net16),
    .C1(net62),
    .D1(net947),
    .Y(net67));
 sky130_fd_sc_hd__a2111o_1 c131 (.A1(net65),
    .A2(net947),
    .B1(net902),
    .C1(net720),
    .D1(net896),
    .X(net68));
 sky130_fd_sc_hd__and3b_2 c132 (.A_N(net818),
    .B(net865),
    .C(net869),
    .X(net69));
 sky130_fd_sc_hd__nor2_4 c133 (.A(net69),
    .B(net811),
    .Y(net70));
 sky130_fd_sc_hd__nand2b_2 c134 (.A_N(net820),
    .B(net69),
    .Y(net71));
 sky130_fd_sc_hd__o2111ai_4 c135 (.A1(net832),
    .A2(net843),
    .B1(net70),
    .C1(net854),
    .D1(net811),
    .Y(net72));
 sky130_fd_sc_hd__nor2_1 c136 (.A(net72),
    .B(net70),
    .Y(net73));
 sky130_fd_sc_hd__and2_1 c137 (.A(net73),
    .B(net817),
    .X(net74));
 sky130_fd_sc_hd__nor2_1 c138 (.A(net819),
    .B(net73),
    .Y(net75));
 sky130_fd_sc_hd__nand2_1 c139 (.A(net75),
    .B(net812),
    .Y(net76));
 sky130_fd_sc_hd__nand3_2 c140 (.A(net813),
    .B(net73),
    .C(net817),
    .Y(net77));
 sky130_fd_sc_hd__nand2b_1 c141 (.A_N(net70),
    .B(net74),
    .Y(net78));
 sky130_fd_sc_hd__and2_4 c142 (.A(net74),
    .B(net78),
    .X(net79));
 sky130_fd_sc_hd__nor2b_2 c143 (.A(net815),
    .B_N(net78),
    .Y(net80));
 sky130_fd_sc_hd__and2_1 c144 (.A(net821),
    .B(net80),
    .X(net81));
 sky130_fd_sc_hd__a2111oi_1 c145 (.A1(net78),
    .A2(net74),
    .B1(net75),
    .C1(net70),
    .D1(net71),
    .Y(net874));
 sky130_fd_sc_hd__and2b_1 c146 (.A_N(net76),
    .B(net80),
    .X(net82));
 sky130_fd_sc_hd__or2_2 c147 (.A(net71),
    .B(net82),
    .X(net83));
 sky130_fd_sc_hd__nor2b_4 c148 (.A(net80),
    .B_N(net81),
    .Y(net84));
 sky130_fd_sc_hd__and2_4 c149 (.A(net82),
    .B(net75),
    .X(net890));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net79),
    .A1(net77),
    .A2(net890),
    .A3(net73),
    .S0(net84),
    .S1(net812),
    .X(net85));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net85),
    .A1(net76),
    .A2(net84),
    .A3(net74),
    .S0(net890),
    .S1(net818),
    .X(net86));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net81),
    .A1(net70),
    .A2(net85),
    .A3(net86),
    .S0(net83),
    .S1(net84),
    .X(net87));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net83),
    .A1(net86),
    .A2(net82),
    .A3(net84),
    .S0(net70),
    .S1(net85),
    .X(net88));
 sky130_fd_sc_hd__or3b_4 c154 (.A(net823),
    .B(net812),
    .C_N(net828),
    .X(net89));
 sky130_fd_sc_hd__nand3b_1 c155 (.A_N(net828),
    .B(net84),
    .C(net72),
    .Y(net90));
 sky130_fd_sc_hd__and3_4 c156 (.A(net831),
    .B(net88),
    .C(net869),
    .X(net91));
 sky130_fd_sc_hd__or3_2 c157 (.A(net90),
    .B(net830),
    .C(net834),
    .X(net92));
 sky130_fd_sc_hd__o2111ai_4 c158 (.A1(net830),
    .A2(net69),
    .B1(net826),
    .C1(net842),
    .D1(net91),
    .Y(net93));
 sky130_fd_sc_hd__nor3b_1 c159 (.A(net93),
    .B(net92),
    .C_N(net829),
    .Y(net94));
 sky130_fd_sc_hd__buf_2 c160 (.A(net674),
    .X(net95));
 sky130_fd_sc_hd__and3b_2 c161 (.A_N(net69),
    .B(net84),
    .C(net836),
    .X(net96));
 sky130_fd_sc_hd__and3b_1 c162 (.A_N(net812),
    .B(net828),
    .C(net842),
    .X(net97));
 sky130_fd_sc_hd__nand3b_4 c163 (.A_N(net824),
    .B(net84),
    .C(net91),
    .Y(net916));
 sky130_fd_sc_hd__nand3b_4 c164 (.A_N(net89),
    .B(net91),
    .C(net72),
    .Y(net98));
 sky130_fd_sc_hd__or3_1 c165 (.A(net98),
    .B(net824),
    .C(net830),
    .X(net99));
 sky130_fd_sc_hd__buf_16 c166 (.A(net674),
    .X(net100));
 sky130_fd_sc_hd__inv_4 c167 (.A(net673),
    .Y(net101));
 sky130_fd_sc_hd__and3_1 c168 (.A(net836),
    .B(net840),
    .C(net97),
    .X(net102));
 sky130_fd_sc_hd__a2111o_4 c169 (.A1(net829),
    .A2(net88),
    .B1(net90),
    .C1(net916),
    .D1(net102),
    .X(net103));
 sky130_fd_sc_hd__sdfrbp_2 c170 (.CLK(clknet_4_2_0_clk),
    .D(net88),
    .RESET_B(net91),
    .SCD(net99),
    .SCE(net95),
    .Q(net105),
    .Q_N(net104));
 sky130_fd_sc_hd__nor3_1 c171 (.A(net102),
    .B(net817),
    .C(net842),
    .Y(net106));
 sky130_fd_sc_hd__a2111oi_2 c172 (.A1(net101),
    .A2(net87),
    .B1(net102),
    .C1(net963),
    .D1(net916),
    .Y(net912));
 sky130_fd_sc_hd__o2111ai_4 c173 (.A1(net814),
    .A2(net916),
    .B1(net101),
    .C1(net963),
    .D1(net89),
    .Y(net107));
 sky130_fd_sc_hd__mux4_4 c174 (.A0(net102),
    .A1(net963),
    .A2(net100),
    .A3(net103),
    .S0(net93),
    .S1(net912),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net103),
    .A1(net94),
    .A2(net96),
    .A3(net963),
    .S0(net100),
    .S1(net1027),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 c176 (.A(net716),
    .X(net110));
 sky130_fd_sc_hd__nor2_2 c177 (.A(net817),
    .B(net100),
    .Y(net111));
 sky130_fd_sc_hd__or2b_4 c178 (.A(net0),
    .B_N(net857),
    .X(net112));
 sky130_fd_sc_hd__and2_1 c179 (.A(net864),
    .B(net111),
    .X(net113));
 sky130_fd_sc_hd__and3_1 c180 (.A(net100),
    .B(net91),
    .C(net858),
    .X(net114));
 sky130_fd_sc_hd__and4b_2 c181 (.A_N(net692),
    .B(net842),
    .C(net960),
    .D(net858),
    .X(net115));
 sky130_fd_sc_hd__and3_1 c182 (.A(net114),
    .B(net79),
    .C(net960),
    .X(net116));
 sky130_fd_sc_hd__sdfrbp_2 c183 (.CLK(clknet_4_8_0_clk),
    .D(net107),
    .RESET_B(net1008),
    .SCD(net112),
    .SCE(net960),
    .Q(net118),
    .Q_N(net117));
 sky130_fd_sc_hd__nor3_2 c184 (.A(net115),
    .B(net977),
    .C(net960),
    .Y(net119));
 sky130_fd_sc_hd__nand3_1 c185 (.A(net111),
    .B(net960),
    .C(net119),
    .Y(net120));
 sky130_fd_sc_hd__and2_1 c186 (.A(net77),
    .B(net2),
    .X(net121));
 sky130_fd_sc_hd__nor4_2 c187 (.A(net121),
    .B(net110),
    .C(net91),
    .D(net960),
    .Y(net122));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net91),
    .A1(net118),
    .A2(net850),
    .A3(net977),
    .S0(net936),
    .S1(net107),
    .X(net123));
 sky130_fd_sc_hd__o2111ai_4 c189 (.A1(net936),
    .A2(net826),
    .B1(net112),
    .C1(net976),
    .D1(net960),
    .Y(net124));
 sky130_fd_sc_hd__nand4_1 c190 (.A(net121),
    .B(net937),
    .C(net117),
    .D(net992),
    .Y(net125));
 sky130_fd_sc_hd__mux4_1 c191 (.A0(net125),
    .A1(net932),
    .A2(net116),
    .A3(net115),
    .S0(net112),
    .S1(net121),
    .X(net126));
 sky130_fd_sc_hd__or4_2 c192 (.A(net848),
    .B(net120),
    .C(net976),
    .D(net916),
    .X(net127));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net118),
    .A1(net124),
    .A2(net937),
    .A3(net127),
    .S0(net107),
    .S1(clknet_1_0__leaf_net725),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net116),
    .A1(net127),
    .A2(net115),
    .A3(net125),
    .S0(net960),
    .S1(net117),
    .X(net129));
 sky130_fd_sc_hd__nand4_1 c195 (.A(net115),
    .B(net937),
    .C(clknet_1_0__leaf_net725),
    .D(clknet_1_0__leaf_net726),
    .Y(net130));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net114),
    .A1(net125),
    .A2(clknet_1_0__leaf_net130),
    .A3(net110),
    .S0(net117),
    .S1(clknet_1_0__leaf_net726),
    .X(net131));
 sky130_fd_sc_hd__sdfbbp_1 c197 (.CLK(clknet_4_8_0_clk),
    .D(net127),
    .RESET_B(net112),
    .SCD(net960),
    .SCE(net706),
    .SET_B(net992),
    .Q(net133),
    .Q_N(net132));
 sky130_fd_sc_hd__inv_1 c198 (.A(net701),
    .Y(net134));
 sky130_fd_sc_hd__nand3_4 c199 (.A(net13),
    .B(net133),
    .C(net17),
    .Y(net135));
 sky130_fd_sc_hd__sdfbbn_1 c200 (.CLK_N(clknet_4_10_0_clk),
    .D(net853),
    .RESET_B(net22),
    .SCD(net98),
    .SCE(net857),
    .SET_B(net931),
    .Q(net137),
    .Q_N(net136));
 sky130_fd_sc_hd__or3_2 c201 (.A(net960),
    .B(net706),
    .C(net1027),
    .X(net138));
 sky130_fd_sc_hd__nor3_2 c202 (.A(net84),
    .B(net8),
    .C(net853),
    .Y(net139));
 sky130_fd_sc_hd__nor3b_2 c203 (.A(net139),
    .B(net858),
    .C_N(net25),
    .Y(net140));
 sky130_fd_sc_hd__dlygate4sd1_1 c204 (.A(net701),
    .X(net141));
 sky130_fd_sc_hd__buf_2 c205 (.A(net711),
    .X(net142));
 sky130_fd_sc_hd__inv_4 c206 (.A(net716),
    .Y(net143));
 sky130_fd_sc_hd__nand3b_1 c207 (.A_N(net826),
    .B(net140),
    .C(net1027),
    .Y(net144));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(net18),
    .A1(net143),
    .A2(net144),
    .A3(net976),
    .S0(net142),
    .S1(net141),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net23),
    .A1(net115),
    .A2(net105),
    .A3(net141),
    .S0(net103),
    .S1(net134),
    .X(net146));
 sky130_fd_sc_hd__mux4_4 c210 (.A0(net17),
    .A1(net145),
    .A2(net826),
    .A3(net98),
    .S0(net18),
    .S1(clknet_1_0__leaf_net727),
    .X(net147));
 sky130_fd_sc_hd__nor3_2 c211 (.A(net19),
    .B(net916),
    .C(clknet_1_1__leaf_net727),
    .Y(net148));
 sky130_fd_sc_hd__clkbuf_2 c212 (.A(net700),
    .X(net149));
 sky130_fd_sc_hd__mux4_2 c213 (.A0(net149),
    .A1(net143),
    .A2(net25),
    .A3(net145),
    .S0(net937),
    .S1(net144),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net144),
    .A1(net13),
    .A2(net149),
    .A3(net844),
    .S0(net138),
    .S1(clknet_1_0__leaf_net727),
    .X(net151));
 sky130_fd_sc_hd__or3b_2 c215 (.A(net143),
    .B(clknet_1_0__leaf_net151),
    .C_N(net17),
    .X(net152));
 sky130_fd_sc_hd__a2111o_1 c216 (.A1(clknet_1_1__leaf_net152),
    .A2(clknet_1_0__leaf_net151),
    .B1(net17),
    .C1(net961),
    .D1(net135),
    .X(net153));
 sky130_fd_sc_hd__clkinv_2 c217 (.A(net807),
    .Y(net154));
 sky130_fd_sc_hd__mux4_2 c218 (.A0(net134),
    .A1(clknet_1_0__leaf_net152),
    .A2(clknet_1_1__leaf_net151),
    .A3(net150),
    .S0(net154),
    .S1(net25),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net154),
    .A1(clknet_1_0__leaf_net153),
    .A2(clknet_1_0__leaf_net152),
    .A3(net142),
    .S0(net145),
    .S1(clknet_1_1__leaf_net727),
    .X(net156));
 sky130_fd_sc_hd__or3b_1 c220 (.A(net33),
    .B(net136),
    .C_N(net731),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 c221 (.A(net1019),
    .X(net158));
 sky130_fd_sc_hd__buf_16 c222 (.A(net795),
    .X(net884));
 sky130_fd_sc_hd__nor3_2 c223 (.A(net857),
    .B(net861),
    .C(net138),
    .Y(net159));
 sky130_fd_sc_hd__nor3b_1 c224 (.A(net138),
    .B(net120),
    .C_N(net976),
    .Y(net160));
 sky130_fd_sc_hd__or3b_4 c225 (.A(net950),
    .B(net25),
    .C_N(net729),
    .X(net895));
 sky130_fd_sc_hd__and3_1 c226 (.A(net157),
    .B(net890),
    .C(net37),
    .X(net161));
 sky130_fd_sc_hd__nor2b_1 c227 (.A(net137),
    .B_N(net728),
    .Y(net162));
 sky130_fd_sc_hd__buf_2 c228 (.A(net660),
    .X(net898));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net98),
    .A1(net834),
    .A2(net132),
    .A3(net160),
    .S0(net29),
    .S1(net43),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 c230 (.A(net902),
    .X(net164));
 sky130_fd_sc_hd__nor3_1 c231 (.A(net164),
    .B(net916),
    .C(net898),
    .Y(net165));
 sky130_fd_sc_hd__nand3b_1 c232 (.A_N(net120),
    .B(net149),
    .C(net898),
    .Y(net166));
 sky130_fd_sc_hd__and4bb_1 c233 (.A_N(net161),
    .B_N(net930),
    .C(net19),
    .D(net962),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 c234 (.A(net659),
    .X(net168));
 sky130_fd_sc_hd__or3_4 c235 (.A(net166),
    .B(net98),
    .C(net728),
    .X(net169));
 sky130_fd_sc_hd__dfbbn_1 c236 (.CLK_N(clknet_4_10_0_clk),
    .D(net19),
    .RESET_B(net931),
    .SET_B(net169),
    .Q(net171),
    .Q_N(net170));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net163),
    .A1(net168),
    .A2(net171),
    .A3(net169),
    .S0(net29),
    .S1(net138),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net158),
    .A1(net168),
    .A2(net29),
    .A3(net950),
    .S0(net169),
    .S1(net1009),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net162),
    .A1(net168),
    .A2(net930),
    .A3(net170),
    .S0(net729),
    .S1(net1001),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net884),
    .A1(net29),
    .A2(net895),
    .A3(net687),
    .S0(net715),
    .S1(net733),
    .X(net175));
 sky130_fd_sc_hd__mux4_2 c241 (.A0(net175),
    .A1(net895),
    .A2(net168),
    .A3(net161),
    .S0(net715),
    .S1(net732),
    .X(net918));
 sky130_fd_sc_hd__nand2_1 c242 (.A(net175),
    .B(net50),
    .Y(net176));
 sky130_fd_sc_hd__nor2b_1 c243 (.A(net68),
    .B_N(net896),
    .Y(net177));
 sky130_fd_sc_hd__a2111o_4 c244 (.A1(net46),
    .A2(net68),
    .B1(net50),
    .C1(net962),
    .D1(net54),
    .X(net178));
 sky130_fd_sc_hd__or3_2 c245 (.A(net68),
    .B(net688),
    .C(net721),
    .X(net179));
 sky130_fd_sc_hd__nor2b_1 c246 (.A(net950),
    .B_N(net54),
    .Y(net920));
 sky130_fd_sc_hd__and2b_1 c247 (.A_N(net61),
    .B(net178),
    .X(net180));
 sky130_fd_sc_hd__nand3b_1 c248 (.A_N(net947),
    .B(net179),
    .C(net962),
    .Y(net181));
 sky130_fd_sc_hd__clkbuf_1 c249 (.A(net798),
    .X(net182));
 sky130_fd_sc_hd__sdfbbn_1 c250 (.CLK_N(clknet_4_10_0_clk),
    .D(net178),
    .RESET_B(net861),
    .SCD(net895),
    .SCE(net169),
    .SET_B(net721),
    .Q(net921),
    .Q_N(net183));
 sky130_fd_sc_hd__buf_16 c251 (.A(net798),
    .X(net888));
 sky130_fd_sc_hd__o2111a_1 c252 (.A1(net181),
    .A2(net46),
    .B1(net962),
    .C1(net183),
    .D1(net62),
    .X(net184));
 sky130_fd_sc_hd__nor2b_2 c253 (.A(net52),
    .B_N(net46),
    .Y(net892));
 sky130_fd_sc_hd__a2111oi_1 c254 (.A1(net57),
    .A2(net169),
    .B1(net892),
    .C1(net61),
    .D1(net730),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 c255 (.A(net808),
    .Y(net910));
 sky130_fd_sc_hd__o2111ai_1 c256 (.A1(net62),
    .A2(net55),
    .B1(net178),
    .C1(net891),
    .D1(net56),
    .Y(net186));
 sky130_fd_sc_hd__and2_0 c257 (.A(net1017),
    .B(net731),
    .X(net187));
 sky130_fd_sc_hd__o2111a_1 c258 (.A1(net179),
    .A2(net892),
    .B1(net56),
    .C1(net947),
    .D1(net731),
    .X(net919));
 sky130_fd_sc_hd__or3b_1 c259 (.A(net182),
    .B(net50),
    .C_N(net913),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net188),
    .A1(net183),
    .A2(net947),
    .A3(net68),
    .S0(net178),
    .S1(net54),
    .X(net899));
 sky130_fd_sc_hd__sdfbbp_1 c261 (.CLK(clknet_4_10_0_clk),
    .D(net187),
    .RESET_B(net184),
    .SCD(net899),
    .SCE(net179),
    .SET_B(net947),
    .Q(net917),
    .Q_N(net189));
 sky130_fd_sc_hd__o2111ai_4 c262 (.A1(net176),
    .A2(net189),
    .B1(net921),
    .C1(net178),
    .D1(net52),
    .Y(net909));
 sky130_fd_sc_hd__o2111a_1 c263 (.A1(net177),
    .A2(net909),
    .B1(net189),
    .C1(net57),
    .D1(net861),
    .X(net190));
 sky130_fd_sc_hd__nor3b_1 c264 (.A(net76),
    .B(net818),
    .C_N(net85),
    .Y(net191));
 sky130_fd_sc_hd__or2b_1 c265 (.A(net870),
    .B_N(net1025),
    .X(net192));
 sky130_fd_sc_hd__and2b_4 c266 (.A_N(net820),
    .B(net191),
    .X(net193));
 sky130_fd_sc_hd__and2_1 c267 (.A(net81),
    .B(net70),
    .X(net194));
 sky130_fd_sc_hd__nor2b_1 c268 (.A(net635),
    .B_N(net193),
    .Y(net195));
 sky130_fd_sc_hd__and3b_1 c269 (.A_N(net80),
    .B(net955),
    .C(net85),
    .X(net196));
 sky130_fd_sc_hd__nand2b_1 c270 (.A_N(net193),
    .B(net70),
    .Y(net197));
 sky130_fd_sc_hd__a2111o_1 c271 (.A1(net193),
    .A2(net77),
    .B1(net71),
    .C1(net72),
    .D1(net81),
    .X(net198));
 sky130_fd_sc_hd__or2_1 c272 (.A(net88),
    .B(net76),
    .X(net199));
 sky130_fd_sc_hd__nor2_1 c273 (.A(net198),
    .B(net943),
    .Y(net200));
 sky130_fd_sc_hd__and3_2 c274 (.A(net200),
    .B(net199),
    .C(net194),
    .X(net201));
 sky130_fd_sc_hd__or3b_1 c275 (.A(net196),
    .B(net200),
    .C_N(net943),
    .X(net202));
 sky130_fd_sc_hd__buf_2 c276 (.A(net712),
    .X(net203));
 sky130_fd_sc_hd__or3_1 c277 (.A(net194),
    .B(net198),
    .C(net943),
    .X(net204));
 sky130_fd_sc_hd__a2111o_1 c278 (.A1(net204),
    .A2(net192),
    .B1(net943),
    .C1(net85),
    .D1(net1026),
    .X(net205));
 sky130_fd_sc_hd__o2111a_1 c279 (.A1(net943),
    .A2(net820),
    .B1(net201),
    .C1(net81),
    .D1(net1026),
    .X(net206));
 sky130_fd_sc_hd__sdfrtn_1 c280 (.CLK_N(clknet_4_0_0_clk),
    .D(net205),
    .RESET_B(net194),
    .SCD(net943),
    .SCE(net1026),
    .Q(net207));
 sky130_fd_sc_hd__and3_2 c281 (.A(net204),
    .B(net1026),
    .C(net1003),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net195),
    .A1(net202),
    .A2(net208),
    .A3(net201),
    .S0(net72),
    .S1(net193),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net208),
    .A1(net207),
    .A2(net202),
    .A3(net201),
    .S0(net1026),
    .S1(net681),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net202),
    .A1(net83),
    .A2(net86),
    .A3(net943),
    .S0(net945),
    .S1(net973),
    .X(net211));
 sky130_fd_sc_hd__sdfbbn_1 c285 (.CLK_N(clknet_4_0_0_clk),
    .D(net1000),
    .RESET_B(net208),
    .SCD(net682),
    .SCE(net973),
    .SET_B(net993),
    .Q(net213),
    .Q_N(net212));
 sky130_fd_sc_hd__and2b_1 c286 (.A_N(net196),
    .B(net844),
    .X(net214));
 sky130_fd_sc_hd__nor2_2 c287 (.A(net192),
    .B(net92),
    .Y(net215));
 sky130_fd_sc_hd__nand2b_1 c288 (.A_N(net72),
    .B(net1026),
    .Y(net216));
 sky130_fd_sc_hd__or2_4 c289 (.A(net101),
    .B(net77),
    .X(net217));
 sky130_fd_sc_hd__or2_1 c290 (.A(net195),
    .B(net214),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 c291 (.A(net707),
    .X(net219));
 sky130_fd_sc_hd__o2111a_2 c292 (.A1(net218),
    .A2(net825),
    .B1(net193),
    .C1(net104),
    .D1(net1027),
    .X(net220));
 sky130_fd_sc_hd__or3b_1 c293 (.A(net105),
    .B(net682),
    .C_N(net723),
    .X(net221));
 sky130_fd_sc_hd__and3b_1 c294 (.A_N(net214),
    .B(net219),
    .C(net218),
    .X(net222));
 sky130_fd_sc_hd__or2_1 c295 (.A(net218),
    .B(net196),
    .X(net223));
 sky130_fd_sc_hd__inv_2 c296 (.A(net707),
    .Y(net224));
 sky130_fd_sc_hd__buf_2 c297 (.A(net673),
    .X(net225));
 sky130_fd_sc_hd__buf_6 c298 (.A(net712),
    .X(net226));
 sky130_fd_sc_hd__buf_1 c299 (.A(net806),
    .X(net227));
 sky130_fd_sc_hd__a2111o_2 c300 (.A1(net106),
    .A2(net197),
    .B1(net968),
    .C1(net95),
    .D1(net840),
    .X(net228));
 sky130_fd_sc_hd__a2111oi_1 c301 (.A1(net968),
    .A2(net219),
    .B1(net226),
    .C1(net72),
    .D1(net220),
    .Y(net229));
 sky130_fd_sc_hd__mux4_2 c302 (.A0(net221),
    .A1(net916),
    .A2(net955),
    .A3(net97),
    .S0(net217),
    .S1(net1027),
    .X(net230));
 sky130_fd_sc_hd__inv_6 c303 (.A(net809),
    .Y(net231));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net223),
    .A1(net221),
    .A2(net217),
    .A3(net201),
    .S0(net72),
    .S1(net968),
    .X(net232));
 sky130_fd_sc_hd__a2111o_4 c305 (.A1(net215),
    .A2(net224),
    .B1(net968),
    .C1(net696),
    .D1(net972),
    .X(net233));
 sky130_fd_sc_hd__a2111oi_1 c306 (.A1(net224),
    .A2(net233),
    .B1(net968),
    .C1(net231),
    .D1(net972),
    .Y(net234));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net201),
    .A1(net935),
    .A2(net233),
    .A3(net847),
    .S0(net230),
    .S1(net987),
    .X(net235));
 sky130_fd_sc_hd__or3b_4 c308 (.A(net838),
    .B(net227),
    .C_N(net696),
    .X(net236));
 sky130_fd_sc_hd__buf_4 c309 (.A(clknet_1_0__leaf_net800),
    .X(net237));
 sky130_fd_sc_hd__and4b_1 c310 (.A_N(net865),
    .B(net935),
    .C(net862),
    .D(net236),
    .X(net238));
 sky130_fd_sc_hd__nor4_1 c311 (.A(net110),
    .B(net119),
    .C(net696),
    .D(net724),
    .Y(net239));
 sky130_fd_sc_hd__and2_1 c312 (.A(net239),
    .B(net724),
    .X(net240));
 sky130_fd_sc_hd__o2111a_1 c313 (.A1(net127),
    .A2(net112),
    .B1(net236),
    .C1(net1010),
    .D1(net973),
    .X(net241));
 sky130_fd_sc_hd__or4b_1 c314 (.A(net112),
    .B(net236),
    .C(net110),
    .D_N(net961),
    .X(net242));
 sky130_fd_sc_hd__nor2_1 c315 (.A(net825),
    .B(net215),
    .Y(net243));
 sky130_fd_sc_hd__nand4_2 c316 (.A(net242),
    .B(net240),
    .C(net236),
    .D(net916),
    .Y(net244));
 sky130_fd_sc_hd__or2_2 c317 (.A(net197),
    .B(clknet_1_0__leaf_net726),
    .X(net245));
 sky130_fd_sc_hd__and2b_1 c318 (.A_N(net87),
    .B(net227),
    .X(net246));
 sky130_fd_sc_hd__and3_2 c319 (.A(net240),
    .B(clknet_1_0__leaf_net245),
    .C(net239),
    .X(net247));
 sky130_fd_sc_hd__and4bb_1 c320 (.A_N(net207),
    .B_N(net236),
    .C(net942),
    .D(net112),
    .X(net248));
 sky130_fd_sc_hd__nor4b_1 c321 (.A(net237),
    .B(net231),
    .C(net236),
    .D_N(net942),
    .Y(net249));
 sky130_fd_sc_hd__sdfrtp_4 c322 (.CLK(clknet_4_2_0_clk),
    .D(net119),
    .RESET_B(net238),
    .SCD(clknet_1_0__leaf_net247),
    .SCE(net231),
    .Q(net250));
 sky130_fd_sc_hd__mux4_2 c323 (.A0(net248),
    .A1(net942),
    .A2(net825),
    .A3(net858),
    .S0(net862),
    .S1(net987),
    .X(net251));
 sky130_fd_sc_hd__nor4_1 c324 (.A(net227),
    .B(net250),
    .C(clknet_1_0__leaf_net245),
    .D(net217),
    .Y(net252));
 sky130_fd_sc_hd__sdfrtp_1 c325 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_1__leaf_net249),
    .RESET_B(net112),
    .SCD(clknet_1_1__leaf_net252),
    .SCE(net929),
    .Q(net253));
 sky130_fd_sc_hd__sdfrtp_2 c326 (.CLK(clknet_4_2_0_clk),
    .D(net238),
    .RESET_B(net991),
    .SCD(clknet_1_0__leaf_net247),
    .SCE(clknet_1_0__leaf_net249),
    .Q(net254));
 sky130_fd_sc_hd__a2111oi_1 c327 (.A1(net92),
    .A2(clknet_1_1__leaf_net247),
    .B1(net251),
    .C1(net254),
    .D1(net253),
    .Y(net255));
 sky130_fd_sc_hd__sdfbbn_1 c328 (.CLK_N(clknet_4_3_0_clk),
    .D(net929),
    .RESET_B(net243),
    .SCD(net254),
    .SCE(clknet_1_0__leaf_net252),
    .SET_B(net923),
    .Q(net257),
    .Q_N(net256));
 sky130_fd_sc_hd__mux4_2 c329 (.A0(net251),
    .A1(net253),
    .A2(net254),
    .A3(clknet_1_1__leaf_net252),
    .S0(net929),
    .S1(net923),
    .X(net258));
 sky130_fd_sc_hd__or3_1 c330 (.A(net154),
    .B(net141),
    .C(net140),
    .X(net259));
 sky130_fd_sc_hd__or3b_1 c331 (.A(net122),
    .B(net217),
    .C_N(net141),
    .X(net260));
 sky130_fd_sc_hd__and3_1 c332 (.A(clknet_1_1__leaf_net152),
    .B(net203),
    .C(net887),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 c333 (.A(net711),
    .X(net262));
 sky130_fd_sc_hd__buf_8 c334 (.A(net711),
    .X(net881));
 sky130_fd_sc_hd__and3b_2 c335 (.A_N(net141),
    .B(net961),
    .C(net923),
    .X(net903));
 sky130_fd_sc_hd__buf_2 c336 (.A(net805),
    .X(net263));
 sky130_fd_sc_hd__nor3b_1 c337 (.A(net253),
    .B(net263),
    .C_N(net942),
    .Y(net264));
 sky130_fd_sc_hd__mux4_2 c338 (.A0(net148),
    .A1(net263),
    .A2(net890),
    .A3(net881),
    .S0(net259),
    .S1(net961),
    .X(net265));
 sky130_fd_sc_hd__mux4_4 c339 (.A0(net263),
    .A1(net977),
    .A2(net929),
    .A3(net956),
    .S0(net22),
    .S1(net260),
    .X(net266));
 sky130_fd_sc_hd__o2111a_1 c340 (.A1(net263),
    .A2(net881),
    .B1(net104),
    .C1(net699),
    .D1(net736),
    .X(net267));
 sky130_fd_sc_hd__nand3b_4 c341 (.A_N(net142),
    .B(net263),
    .C(net736),
    .Y(net871));
 sky130_fd_sc_hd__or3b_1 c342 (.A(net263),
    .B(net976),
    .C_N(net736),
    .X(net268));
 sky130_fd_sc_hd__mux4_4 c343 (.A0(net268),
    .A1(net122),
    .A2(net150),
    .A3(net135),
    .S0(net5),
    .S1(net267),
    .X(net269));
 sky130_fd_sc_hd__o2111a_4 c344 (.A1(clknet_1_1__leaf_net153),
    .A2(net268),
    .B1(net263),
    .C1(net871),
    .D1(net736),
    .X(net270));
 sky130_fd_sc_hd__or3_4 c345 (.A(net264),
    .B(net262),
    .C(net738),
    .X(net271));
 sky130_fd_sc_hd__sdfbbp_1 c346 (.CLK(clknet_4_8_0_clk),
    .D(net267),
    .RESET_B(net4),
    .SCD(net271),
    .SCE(net103),
    .SET_B(net998),
    .Q(net273),
    .Q_N(net272));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net273),
    .A1(clknet_1_0__leaf_net261),
    .A2(net79),
    .A3(net264),
    .S0(net699),
    .S1(net736),
    .X(net274));
 sky130_fd_sc_hd__inv_6 c348 (.A(net711),
    .Y(net275));
 sky130_fd_sc_hd__o2111a_1 c349 (.A1(net275),
    .A2(net137),
    .B1(net154),
    .C1(net871),
    .D1(net737),
    .X(net276));
 sky130_fd_sc_hd__mux4_4 c350 (.A0(net273),
    .A1(net275),
    .A2(net871),
    .A3(net271),
    .S0(net699),
    .S1(net738),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net262),
    .A1(net264),
    .A2(net275),
    .A3(net271),
    .S0(net737),
    .S1(net1014),
    .X(net278));
 sky130_fd_sc_hd__inv_1 c352 (.A(net797),
    .Y(net279));
 sky130_fd_sc_hd__clkbuf_1 c353 (.A(net797),
    .X(net280));
 sky130_fd_sc_hd__sdfsbp_1 c354 (.CLK(clknet_4_11_0_clk),
    .D(net930),
    .SCD(net25),
    .SCE(net42),
    .SET_B(net159),
    .Q(net282),
    .Q_N(net281));
 sky130_fd_sc_hd__nor4_1 c355 (.A(net279),
    .B(net118),
    .C(net891),
    .D(net271),
    .Y(net283));
 sky130_fd_sc_hd__or4b_2 c356 (.A(net280),
    .B(net942),
    .C(net250),
    .D_N(net987),
    .X(net284));
 sky130_fd_sc_hd__nand4b_4 c357 (.A_N(net282),
    .B(net31),
    .C(net293),
    .D(net887),
    .Y(net285));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net29),
    .A1(net279),
    .A2(net284),
    .A3(net285),
    .S0(net956),
    .S1(net43),
    .X(net286));
 sky130_fd_sc_hd__buf_6 c359 (.A(net799),
    .X(net873));
 sky130_fd_sc_hd__sdfbbn_2 c360 (.CLK_N(clknet_4_11_0_clk),
    .D(net293),
    .RESET_B(net873),
    .SCD(net285),
    .SCE(net890),
    .SET_B(net169),
    .Q(net288),
    .Q_N(net287));
 sky130_fd_sc_hd__inv_2 c361 (.A(net700),
    .Y(net289));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net271),
    .A1(net884),
    .A2(net916),
    .A3(net281),
    .S0(net956),
    .S1(net170),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net295),
    .A1(net282),
    .A2(net288),
    .A3(net873),
    .S0(net25),
    .S1(net907),
    .X(net291));
 sky130_fd_sc_hd__and3_2 c364 (.A(net873),
    .B(net291),
    .C(net742),
    .X(net885));
 sky130_fd_sc_hd__mux4_2 c365 (.A0(net291),
    .A1(net956),
    .A2(net873),
    .A3(net285),
    .S0(net885),
    .S1(net907),
    .X(net292));
 sky130_fd_sc_hd__mux4_2 c366 (.A0(net171),
    .A1(net288),
    .A2(net873),
    .A3(net236),
    .S0(net289),
    .S1(net688),
    .X(net878));
 sky130_fd_sc_hd__and3b_1 c367 (.A_N(net25),
    .B(net871),
    .C(net170),
    .X(net293));
 sky130_fd_sc_hd__inv_2 c368 (.A(net799),
    .Y(net294));
 sky130_fd_sc_hd__nor3_1 c369 (.A(net39),
    .B(net41),
    .C(net25),
    .Y(net295));
 sky130_fd_sc_hd__mux4_2 c370 (.A0(net289),
    .A1(net950),
    .A2(net39),
    .A3(net885),
    .S0(net834),
    .S1(net878),
    .X(net900));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net288),
    .A1(net863),
    .A2(net885),
    .A3(net962),
    .S0(net950),
    .S1(net742),
    .X(net296));
 sky130_fd_sc_hd__mux4_2 c372 (.A0(net294),
    .A1(net834),
    .A2(net289),
    .A3(net838),
    .S0(net292),
    .S1(net900),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net286),
    .A1(net296),
    .A2(net900),
    .A3(net297),
    .S0(net847),
    .S1(net31),
    .X(net298));
 sky130_fd_sc_hd__mux4_4 c392 (.A0(net169),
    .A1(net909),
    .A2(net881),
    .A3(net892),
    .S0(net915),
    .S1(net907),
    .X(net299));
 sky130_fd_sc_hd__mux4_2 c393 (.A0(net276),
    .A1(net240),
    .A2(net962),
    .A3(net909),
    .S0(net61),
    .S1(clknet_1_0__leaf_net908),
    .X(net300));
 sky130_fd_sc_hd__mux4_4 c394 (.A0(net157),
    .A1(net899),
    .A2(net891),
    .A3(net913),
    .S1(clknet_1_0__leaf_net908),
    .X(net301));
 sky130_fd_sc_hd__a2111o_1 c395 (.A1(net962),
    .A2(net61),
    .B1(net917),
    .C1(net925),
    .D1(clknet_1_1__leaf_net908),
    .X(net897));
 sky130_fd_sc_hd__nor2b_2 c396 (.A(net70),
    .B_N(net735),
    .Y(net302));
 sky130_fd_sc_hd__clkbuf_2 c397 (.A(net1007),
    .X(net303));
 sky130_fd_sc_hd__nand2b_1 c398 (.A_N(net303),
    .B(net819),
    .Y(net304));
 sky130_fd_sc_hd__and3b_1 c399 (.A_N(net943),
    .B(net869),
    .C(net198),
    .X(net305));
 sky130_fd_sc_hd__or2b_2 c400 (.A(net85),
    .B_N(net199),
    .X(net306));
 sky130_fd_sc_hd__nor2_2 c401 (.A(net305),
    .B(net85),
    .Y(net307));
 sky130_fd_sc_hd__nand2b_2 c402 (.A_N(net305),
    .B(net306),
    .Y(net308));
 sky130_fd_sc_hd__inv_1 c403 (.A(net676),
    .Y(net309));
 sky130_fd_sc_hd__inv_6 c404 (.A(net663),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 c405 (.A(net663),
    .Y(net311));
 sky130_fd_sc_hd__and2_1 c406 (.A(net310),
    .B(net311),
    .X(net312));
 sky130_fd_sc_hd__or2_1 c407 (.A(net945),
    .B(net303),
    .X(net313));
 sky130_fd_sc_hd__nor4_1 c408 (.A(net309),
    .B(net312),
    .C(net310),
    .D(net944),
    .Y(net314));
 sky130_fd_sc_hd__mux4_1 c409 (.A0(net304),
    .A1(net302),
    .A2(net312),
    .A3(net307),
    .S0(net309),
    .S1(net310),
    .X(net315));
 sky130_fd_sc_hd__o2111ai_2 c410 (.A1(net311),
    .A2(net302),
    .B1(net1026),
    .C1(net735),
    .D1(clknet_1_0__leaf_net743),
    .Y(net316));
 sky130_fd_sc_hd__or2_2 c411 (.A(net303),
    .B(clknet_1_0__leaf_net743),
    .X(net317));
 sky130_fd_sc_hd__sdfsbp_1 c412 (.CLK(clknet_4_1_0_clk),
    .D(net306),
    .SCD(net308),
    .SCE(net943),
    .SET_B(net193),
    .Q(net319),
    .Q_N(net318));
 sky130_fd_sc_hd__mux4_4 c413 (.A0(net944),
    .A1(clknet_1_0__leaf_net316),
    .A2(net319),
    .A3(net308),
    .S0(net939),
    .S1(net311),
    .X(net320));
 sky130_fd_sc_hd__mux4_4 c414 (.A0(clknet_1_0__leaf_net317),
    .A1(net944),
    .A2(net307),
    .A3(net312),
    .S0(net939),
    .S1(clknet_1_0__leaf_net744),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net306),
    .A1(clknet_1_1__leaf_net317),
    .A2(net944),
    .A3(net939),
    .S0(clknet_1_0__leaf_net744),
    .S1(net746),
    .X(net322));
 sky130_fd_sc_hd__mux4_4 c416 (.A0(clknet_1_1__leaf_net316),
    .A1(net318),
    .A2(net312),
    .A3(clknet_1_0__leaf_net322),
    .S0(clknet_1_0__leaf_net744),
    .S1(net745),
    .X(net323));
 sky130_fd_sc_hd__sdfbbn_1 c417 (.CLK_N(clknet_4_1_0_clk),
    .D(net312),
    .RESET_B(clknet_1_0__leaf_net322),
    .SCD(net85),
    .SCE(net939),
    .SET_B(net746),
    .Q(net325),
    .Q_N(net324));
 sky130_fd_sc_hd__clkbuf_1 c418 (.A(net631),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 c419 (.A(net631),
    .X(net327));
 sky130_fd_sc_hd__nor2b_1 c420 (.A(net869),
    .B_N(net233),
    .Y(net328));
 sky130_fd_sc_hd__nor2b_1 c421 (.A(net95),
    .B_N(net818),
    .Y(net329));
 sky130_fd_sc_hd__clkbuf_1 c422 (.A(net714),
    .X(net330));
 sky130_fd_sc_hd__buf_8 c423 (.A(net809),
    .X(net331));
 sky130_fd_sc_hd__and3_4 c424 (.A(net972),
    .B(net331),
    .C(net304),
    .X(net332));
 sky130_fd_sc_hd__or4b_1 c425 (.A(net327),
    .B(net222),
    .C(net1026),
    .D_N(net1007),
    .X(net333));
 sky130_fd_sc_hd__inv_2 c426 (.A(net713),
    .Y(net334));
 sky130_fd_sc_hd__or3_4 c427 (.A(net1027),
    .B(net332),
    .C(net1026),
    .X(net335));
 sky130_fd_sc_hd__or3_4 c428 (.A(net312),
    .B(net326),
    .C(net335),
    .X(net336));
 sky130_fd_sc_hd__or2_4 c429 (.A(net309),
    .B(net332),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net334),
    .A1(net331),
    .A2(net934),
    .A3(net587),
    .S0(net79),
    .S1(net723),
    .X(net338));
 sky130_fd_sc_hd__inv_1 c431 (.A(net714),
    .Y(net339));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net338),
    .A1(net95),
    .A2(net337),
    .A3(net329),
    .S0(net1027),
    .S1(clknet_1_0__leaf_net743),
    .X(net340));
 sky130_fd_sc_hd__nand3_4 c433 (.A(net336),
    .B(net331),
    .C(net972),
    .Y(net341));
 sky130_fd_sc_hd__nor3_1 c434 (.A(net329),
    .B(net324),
    .C(net336),
    .Y(net342));
 sky130_fd_sc_hd__or2b_1 c435 (.A(net339),
    .B_N(net332),
    .X(net343));
 sky130_fd_sc_hd__a2111oi_2 c436 (.A1(net342),
    .A2(net335),
    .B1(net309),
    .C1(net337),
    .D1(net685),
    .Y(net344));
 sky130_fd_sc_hd__and3_1 c437 (.A(net327),
    .B(net344),
    .C(net1026),
    .X(net345));
 sky130_fd_sc_hd__mux4_2 c438 (.A0(net345),
    .A1(net331),
    .A2(net342),
    .A3(net363),
    .S0(net327),
    .S1(net104),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net344),
    .A1(net346),
    .A2(net337),
    .A3(net220),
    .S0(net834),
    .S1(net684),
    .X(net347));
 sky130_fd_sc_hd__nand2_1 c440 (.A(net325),
    .B(net1005),
    .Y(net348));
 sky130_fd_sc_hd__inv_4 c441 (.A(net712),
    .Y(net349));
 sky130_fd_sc_hd__and4b_4 c442 (.A_N(net243),
    .B(net325),
    .C(net331),
    .D(clknet_1_0__leaf_net726),
    .X(net350));
 sky130_fd_sc_hd__sdfstp_2 c443 (.CLK(clknet_4_9_0_clk),
    .D(net929),
    .SCD(net337),
    .SCE(clknet_1_0__leaf_net252),
    .SET_B(net992),
    .Q(net351));
 sky130_fd_sc_hd__and4_1 c444 (.A(net348),
    .B(net335),
    .C(net341),
    .D(net887),
    .X(net352));
 sky130_fd_sc_hd__buf_6 c445 (.A(net640),
    .X(net353));
 sky130_fd_sc_hd__or2b_2 c446 (.A(net226),
    .B_N(net303),
    .X(net354));
 sky130_fd_sc_hd__nor4_4 c447 (.A(clknet_1_0__leaf_net350),
    .B(net351),
    .C(net353),
    .D(clknet_1_1__leaf_net725),
    .Y(net355));
 sky130_fd_sc_hd__nor2b_1 c448 (.A(net352),
    .B_N(net734),
    .Y(net356));
 sky130_fd_sc_hd__nand4_1 c449 (.A(net840),
    .B(net942),
    .C(net348),
    .D(net203),
    .Y(net357));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net357),
    .A1(net243),
    .A2(net346),
    .A3(net348),
    .S0(net111),
    .S1(net887),
    .X(net358));
 sky130_fd_sc_hd__or2b_2 c451 (.A(net356),
    .B_N(net970),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_2 c452 (.A(net639),
    .X(net360));
 sky130_fd_sc_hd__or2_1 c453 (.A(net346),
    .B(net939),
    .X(net361));
 sky130_fd_sc_hd__sdfstp_2 c454 (.CLK(clknet_4_3_0_clk),
    .D(net303),
    .SCD(clknet_1_0__leaf_net355),
    .SCE(net1027),
    .SET_B(clknet_1_1__leaf_net725),
    .Q(net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__sdfbbp_1 c456 (.CLK(clknet_4_3_0_clk),
    .D(net358),
    .RESET_B(net361),
    .SCD(net351),
    .SCE(net357),
    .SET_B(net973),
    .Q(net365),
    .Q_N(net364));
 sky130_fd_sc_hd__mux4_2 c457 (.A0(net344),
    .A1(net365),
    .A2(net844),
    .A3(net362),
    .S0(net226),
    .S1(net337),
    .X(net924));
 sky130_fd_sc_hd__or4_2 c458 (.A(net222),
    .B(net359),
    .C(net360),
    .D(clknet_1_1__leaf_net726),
    .X(net366));
 sky130_fd_sc_hd__or2b_2 c459 (.A(net351),
    .B_N(net879),
    .X(net367));
 sky130_fd_sc_hd__mux4_4 c460 (.A0(net934),
    .A1(net367),
    .A2(net346),
    .A3(net251),
    .S0(net351),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net367),
    .A1(clknet_1_0__leaf_net252),
    .A2(net362),
    .A3(net364),
    .S0(net356),
    .S1(net879),
    .X(net369));
 sky130_fd_sc_hd__buf_4 c462 (.A(clknet_1_0__leaf_net802),
    .X(net370));
 sky130_fd_sc_hd__or3b_4 c463 (.A(net354),
    .B(net341),
    .C_N(clknet_1_1__leaf_net744),
    .X(net371));
 sky130_fd_sc_hd__or3_2 c464 (.A(clknet_1_0__leaf_net370),
    .B(clknet_1_1__leaf_net743),
    .C(clknet_1_1__leaf_net744),
    .X(net372));
 sky130_fd_sc_hd__and3b_1 c465 (.A_N(net361),
    .B(net226),
    .C(net970),
    .X(net373));
 sky130_fd_sc_hd__and3_4 c466 (.A(clknet_1_0__leaf_net370),
    .B(net361),
    .C(net587),
    .X(net374));
 sky130_fd_sc_hd__o2111a_4 c467 (.A1(net374),
    .A2(net135),
    .B1(net942),
    .C1(net861),
    .D1(net203),
    .X(net375));
 sky130_fd_sc_hd__and4b_2 c468 (.A_N(clknet_1_0__leaf_net371),
    .B(clknet_1_0__leaf_net372),
    .C(net970),
    .D(net1027),
    .X(net376));
 sky130_fd_sc_hd__sdfstp_1 c469 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_1__leaf_net372),
    .SCD(clknet_1_0__leaf_net261),
    .SCE(net132),
    .SET_B(net1015),
    .Q(net377));
 sky130_fd_sc_hd__nor4b_2 c470 (.A(clknet_1_1__leaf_net355),
    .B(net354),
    .C(net377),
    .D_N(net337),
    .Y(net378));
 sky130_fd_sc_hd__sedfxbp_1 c471 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net247),
    .DE(net135),
    .SCD(net1016),
    .SCE(clknet_1_1__leaf_net744),
    .Q(net380),
    .Q_N(net379));
 sky130_fd_sc_hd__o2111ai_2 c472 (.A1(net2),
    .A2(clknet_1_1__leaf_net370),
    .B1(net4),
    .C1(net975),
    .D1(net749),
    .Y(net381));
 sky130_fd_sc_hd__o2111ai_1 c473 (.A1(net377),
    .A2(net379),
    .B1(clknet_1_0__leaf_net381),
    .C1(net135),
    .D1(net975),
    .Y(net382));
 sky130_fd_sc_hd__mux4_4 c474 (.A0(net587),
    .A1(clknet_1_0__leaf_net371),
    .A2(net22),
    .A3(net890),
    .S0(clknet_1_0__leaf_net382),
    .S1(clknet_1_0__leaf_net261),
    .X(net383));
 sky130_fd_sc_hd__nor3_4 c475 (.A(net741),
    .B(clknet_1_1__leaf_net381),
    .C(clknet_1_1__leaf_net371),
    .Y(net911));
 sky130_fd_sc_hd__and3_1 c476 (.A(net135),
    .B(net377),
    .C(net79),
    .X(net384));
 sky130_fd_sc_hd__o2111ai_1 c477 (.A1(net236),
    .A2(clknet_1_0__leaf_net381),
    .B1(net5),
    .C1(clknet_1_1__leaf_net371),
    .D1(net750),
    .Y(net385));
 sky130_fd_sc_hd__mux4_2 c478 (.A0(clknet_1_0__leaf_net382),
    .A1(net203),
    .A2(clknet_1_0__leaf_net381),
    .A3(net678),
    .S0(net748),
    .S1(net750),
    .X(net386));
 sky130_fd_sc_hd__a2111oi_2 c479 (.A1(net384),
    .A2(clknet_1_0__leaf_net385),
    .B1(net135),
    .C1(net741),
    .D1(clknet_1_1__leaf_net744),
    .Y(net901));
 sky130_fd_sc_hd__o2111a_2 c480 (.A1(net376),
    .A2(clknet_1_0__leaf_net901),
    .B1(net939),
    .C1(net335),
    .D1(net1027),
    .X(net387));
 sky130_fd_sc_hd__mux4_4 c481 (.A0(net387),
    .A1(net858),
    .A2(clknet_1_0__leaf_net901),
    .A3(net818),
    .S0(net678),
    .S1(net737),
    .X(net906));
 sky130_fd_sc_hd__a2111oi_0 c482 (.A1(clknet_1_0__leaf_net901),
    .A2(net924),
    .B1(net587),
    .C1(net377),
    .D1(net738),
    .Y(net388));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(clknet_1_1__leaf_net385),
    .A1(net388),
    .A2(clknet_1_0__leaf_net382),
    .A3(clknet_1_0__leaf_net906),
    .S0(net881),
    .S1(clknet_1_0__leaf_net901),
    .X(net389));
 sky130_fd_sc_hd__mux4_2 c484 (.A0(net861),
    .A1(net337),
    .A2(net297),
    .A3(net292),
    .S0(net956),
    .S1(net37),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net881),
    .A1(net390),
    .A2(net236),
    .A3(net104),
    .S0(net987),
    .S1(clknet_1_1__leaf_net743),
    .X(net391));
 sky130_fd_sc_hd__mux4_4 c486 (.A0(net133),
    .A1(net43),
    .A2(net285),
    .A3(net168),
    .S0(net390),
    .S1(net22),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net337),
    .A1(net885),
    .A2(net843),
    .A3(net390),
    .S0(net987),
    .S1(net997),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net284),
    .A1(net390),
    .A2(net5),
    .A3(net956),
    .S0(net861),
    .S1(net894),
    .X(net394));
 sky130_fd_sc_hd__mux4_4 c489 (.A0(net171),
    .A1(net390),
    .A2(net895),
    .A3(net985),
    .S0(net354),
    .S1(net971),
    .X(net395));
 sky130_fd_sc_hd__mux4_2 c490 (.A0(net292),
    .A1(net949),
    .A2(net884),
    .A3(net952),
    .S0(net751),
    .S1(net971),
    .X(net396));
 sky130_fd_sc_hd__mux4_2 c491 (.A0(net396),
    .A1(net37),
    .A2(net43),
    .A3(clknet_1_1__leaf_net901),
    .S0(net881),
    .S1(net898),
    .X(net893));
 sky130_fd_sc_hd__mux4_2 c492 (.A0(net168),
    .A1(net133),
    .A2(net881),
    .A3(clknet_1_0__leaf_net911),
    .S0(net118),
    .S1(net753),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net31),
    .A1(net396),
    .A2(net133),
    .A3(net292),
    .S0(net159),
    .S1(net753),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net297),
    .A1(net284),
    .A2(net885),
    .A3(net287),
    .S0(net675),
    .S1(net753),
    .X(net399));
 sky130_fd_sc_hd__mux4_4 c495 (.A0(net159),
    .A1(net285),
    .A2(clknet_1_1__leaf_net381),
    .A3(net396),
    .S0(net390),
    .S1(net753),
    .X(net400));
 sky130_fd_sc_hd__mux4_4 c496 (.A0(net354),
    .A1(net399),
    .A2(net142),
    .A3(clknet_1_1__leaf_net386),
    .S0(net898),
    .S1(net971),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net373),
    .A1(net396),
    .A2(net968),
    .A3(net132),
    .S0(net956),
    .S1(net872),
    .X(net402));
 sky130_fd_sc_hd__mux4_4 c498 (.A0(net142),
    .A1(net292),
    .A2(net337),
    .A3(clknet_1_1__leaf_net386),
    .S0(net871),
    .S1(net971),
    .X(net403));
 sky130_fd_sc_hd__mux4_4 c499 (.A0(net871),
    .A1(net956),
    .A2(net396),
    .A3(net31),
    .S0(clknet_1_1__leaf_net704),
    .S1(net971),
    .X(net880));
 sky130_fd_sc_hd__mux4_2 c500 (.A0(net398),
    .A1(clknet_1_0__leaf_net147),
    .A2(clknet_1_1__leaf_net880),
    .A3(net891),
    .S0(clknet_1_0__leaf_net893),
    .S1(net297),
    .X(net404));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(net217),
    .A1(net390),
    .A2(net398),
    .A3(clknet_1_0__leaf_net901),
    .S0(clknet_1_0__leaf_net880),
    .S1(net754),
    .X(net405));
 sky130_fd_sc_hd__mux4_4 c502 (.A0(net984),
    .A1(clknet_1_1__leaf_net880),
    .A2(net396),
    .A3(net31),
    .S0(net971),
    .S1(net756),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net285),
    .A1(net900),
    .A2(clknet_1_1__leaf_net880),
    .A3(net898),
    .S0(net971),
    .S1(net886),
    .X(net407));
 sky130_fd_sc_hd__o2111a_1 c504 (.A1(clknet_1_0__leaf_net403),
    .A2(clknet_1_0__leaf_net880),
    .B1(net717),
    .C1(net971),
    .D1(net886),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(clknet_1_1__leaf_net403),
    .A1(net895),
    .A2(clknet_1_0__leaf_net704),
    .A3(net753),
    .S0(net755),
    .S1(net886),
    .X(net409));
 sky130_fd_sc_hd__nand3_1 c528 (.A(net213),
    .B(net973),
    .C(net746),
    .Y(net410));
 sky130_fd_sc_hd__nand2_1 c529 (.A(net817),
    .B(net302),
    .Y(net411));
 sky130_fd_sc_hd__a2111o_1 c530 (.A1(net410),
    .A2(net843),
    .B1(net319),
    .C1(net307),
    .D1(net959),
    .X(net412));
 sky130_fd_sc_hd__nor2_4 c531 (.A(net944),
    .B(net735),
    .Y(net413));
 sky130_fd_sc_hd__nand2b_1 c532 (.A_N(net959),
    .B(net697),
    .Y(net414));
 sky130_fd_sc_hd__and2b_2 c533 (.A_N(net86),
    .B(net697),
    .X(net415));
 sky130_fd_sc_hd__or2b_1 c534 (.A(net213),
    .B_N(net939),
    .X(net416));
 sky130_fd_sc_hd__and2b_1 c535 (.A_N(net319),
    .B(net959),
    .X(net417));
 sky130_fd_sc_hd__nor2_1 c536 (.A(net413),
    .B(net818),
    .Y(net418));
 sky130_fd_sc_hd__nor2_2 c537 (.A(net418),
    .B(net939),
    .Y(net419));
 sky130_fd_sc_hd__nor3_1 c538 (.A(net306),
    .B(net417),
    .C(net413),
    .Y(net420));
 sky130_fd_sc_hd__inv_6 c539 (.Y(net421));
 sky130_fd_sc_hd__clkbuf_1 c540 (.A(net636),
    .X(net422));
 sky130_fd_sc_hd__or3b_1 c541 (.A(net421),
    .B(net418),
    .C_N(net302),
    .X(net423));
 sky130_fd_sc_hd__nand2b_1 c542 (.A_N(net416),
    .B(net421),
    .Y(net424));
 sky130_fd_sc_hd__nor4b_1 c543 (.A(net423),
    .B(net212),
    .C(net928),
    .D_N(net413),
    .Y(net425));
 sky130_fd_sc_hd__sedfxbp_2 c544 (.CLK(clknet_4_1_0_clk),
    .D(net424),
    .DE(net421),
    .SCD(net959),
    .SCE(net697),
    .Q(net427),
    .Q_N(net426));
 sky130_fd_sc_hd__nor3b_1 c545 (.A(net426),
    .B(net993),
    .C_N(net745),
    .Y(net428));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net416),
    .A1(net418),
    .A2(net428),
    .A3(net307),
    .S0(net970),
    .S1(net959),
    .X(net429));
 sky130_fd_sc_hd__or3b_2 c547 (.A(net417),
    .B(net416),
    .C_N(net959),
    .X(net430));
 sky130_fd_sc_hd__mux4_4 c548 (.A0(net422),
    .A1(net423),
    .A2(net430),
    .A3(net79),
    .S0(net426),
    .S1(net757),
    .X(net431));
 sky130_fd_sc_hd__mux4_2 c549 (.A0(net418),
    .A1(net416),
    .A2(net318),
    .A3(net970),
    .S0(net697),
    .S1(net757),
    .X(net432));
 sky130_fd_sc_hd__and3b_2 c550 (.A_N(net302),
    .B(net415),
    .C(net747),
    .X(net433));
 sky130_fd_sc_hd__or4b_1 c551 (.A(net427),
    .B(net433),
    .C(net723),
    .D_N(net973),
    .X(net434));
 sky130_fd_sc_hd__nand3_2 c552 (.A(net844),
    .B(net421),
    .C(net427),
    .Y(net435));
 sky130_fd_sc_hd__and3b_2 c553 (.A_N(net421),
    .B(net415),
    .C(net944),
    .X(net436));
 sky130_fd_sc_hd__nor3b_2 c554 (.A(net413),
    .B(net228),
    .C_N(net410),
    .Y(net437));
 sky130_fd_sc_hd__nor3b_4 c555 (.A(net951),
    .B(net944),
    .C_N(net433),
    .Y(net438));
 sky130_fd_sc_hd__and4_1 c556 (.A(net410),
    .B(net421),
    .C(net193),
    .D(net944),
    .X(net439));
 sky130_fd_sc_hd__buf_6 c557 (.A(net693),
    .X(net877));
 sky130_fd_sc_hd__sedfxtp_4 c558 (.CLK(clknet_4_1_0_clk),
    .D(net424),
    .DE(net438),
    .SCD(net944),
    .SCE(net435),
    .Q(net440));
 sky130_fd_sc_hd__and4bb_2 c559 (.A_N(net438),
    .B_N(net427),
    .C(net439),
    .D(net975),
    .X(net441));
 sky130_fd_sc_hd__and4b_1 c560 (.A_N(net439),
    .B(net433),
    .C(net440),
    .D(net313),
    .X(net442));
 sky130_fd_sc_hd__sedfxtp_1 c561 (.CLK(clknet_4_4_0_clk),
    .D(net434),
    .DE(net844),
    .SCD(net441),
    .SCE(net415),
    .Q(net443));
 sky130_fd_sc_hd__mux4_4 c562 (.A0(net417),
    .A1(net443),
    .A2(net437),
    .A3(net440),
    .S0(net434),
    .S1(net413),
    .X(net444));
 sky130_fd_sc_hd__mux4_2 c563 (.A0(net442),
    .A1(net343),
    .A2(net877),
    .A3(net433),
    .S0(net975),
    .S1(net723),
    .X(net445));
 sky130_fd_sc_hd__sdfbbn_1 c564 (.CLK_N(clknet_4_4_0_clk),
    .D(net445),
    .RESET_B(net438),
    .SCD(net440),
    .SCE(net944),
    .SET_B(net427),
    .Q(net447),
    .Q_N(net446));
 sky130_fd_sc_hd__sdfbbn_1 c565 (.CLK_N(clknet_4_4_0_clk),
    .D(net440),
    .RESET_B(net1011),
    .SCD(net1002),
    .SCE(net445),
    .SET_B(net435),
    .Q(net449),
    .Q_N(net448));
 sky130_fd_sc_hd__a2111oi_4 c566 (.A1(net951),
    .A2(net447),
    .B1(net413),
    .C1(net448),
    .D1(clknet_1_0__leaf_net759),
    .Y(net450));
 sky130_fd_sc_hd__mux4_4 c567 (.A0(net193),
    .A1(net445),
    .A2(net443),
    .A3(net446),
    .S0(net415),
    .S1(net426),
    .X(net451));
 sky130_fd_sc_hd__o2111ai_1 c568 (.A1(net443),
    .A2(net441),
    .B1(net445),
    .C1(net449),
    .D1(clknet_1_0__leaf_net759),
    .Y(net452));
 sky130_fd_sc_hd__o2111ai_2 c569 (.A1(net449),
    .A2(net440),
    .B1(net939),
    .C1(net748),
    .D1(clknet_1_0__leaf_net759),
    .Y(net453));
 sky130_fd_sc_hd__mux4_2 c570 (.A0(net447),
    .A1(net877),
    .A2(net193),
    .A3(net951),
    .S0(net442),
    .S1(net694),
    .X(net454));
 sky130_fd_sc_hd__mux4_2 c571 (.A0(net230),
    .A1(clknet_1_0__leaf_net453),
    .A2(net446),
    .A3(net694),
    .S0(clknet_1_0__leaf_net759),
    .S1(clknet_1_0__leaf_net760),
    .X(net455));
 sky130_fd_sc_hd__o2111ai_1 c572 (.A1(net877),
    .A2(net331),
    .B1(net415),
    .C1(net244),
    .D1(clknet_1_1__leaf_net726),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 c573 (.A(net643),
    .Y(net457));
 sky130_fd_sc_hd__or2b_2 c574 (.A(net457),
    .B_N(net349),
    .X(net458));
 sky130_fd_sc_hd__nand3_4 c575 (.A(net331),
    .B(net941),
    .C(clknet_1_1__leaf_net726),
    .Y(net459));
 sky130_fd_sc_hd__a2111o_1 c576 (.A1(net349),
    .A2(net928),
    .B1(net970),
    .C1(net2),
    .D1(net415),
    .X(net460));
 sky130_fd_sc_hd__nor3b_1 c577 (.A(net360),
    .B(net458),
    .C_N(net677),
    .Y(net461));
 sky130_fd_sc_hd__clkbuf_2 c578 (.A(net644),
    .X(net462));
 sky130_fd_sc_hd__nand3b_1 c579 (.A_N(net257),
    .B(net457),
    .C(net359),
    .Y(net463));
 sky130_fd_sc_hd__or4b_4 c580 (.A(net877),
    .B(net462),
    .C(net677),
    .D_N(clknet_1_1__leaf_net760),
    .X(net464));
 sky130_fd_sc_hd__and3_2 c581 (.A(net352),
    .B(net353),
    .C(clknet_1_1__leaf_net726),
    .X(net465));
 sky130_fd_sc_hd__and3b_1 c582 (.A_N(net463),
    .B(net458),
    .C(net433),
    .X(net466));
 sky130_fd_sc_hd__buf_4 c583 (.A(clknet_1_0__leaf_net801),
    .X(net467));
 sky130_fd_sc_hd__nand2b_4 c584 (.A_N(net365),
    .B(clknet_1_0__leaf_net465),
    .Y(net468));
 sky130_fd_sc_hd__nor3b_1 c585 (.A(net458),
    .B(net257),
    .C_N(net747),
    .Y(net469));
 sky130_fd_sc_hd__nor3_1 c586 (.A(net427),
    .B(net970),
    .C(clknet_1_0__leaf_net760),
    .Y(net922));
 sky130_fd_sc_hd__and3_1 c587 (.A(net466),
    .B(net349),
    .C(clknet_1_1__leaf_net760),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 c588 (.A(clknet_1_1__leaf_net800),
    .X(net471));
 sky130_fd_sc_hd__and2_4 c589 (.A(net862),
    .B(clknet_1_1__leaf_net759),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net472),
    .A1(net970),
    .A2(net359),
    .A3(net426),
    .S0(net747),
    .S1(clknet_1_1__leaf_net759),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(clknet_1_1__leaf_net471),
    .A1(net469),
    .A2(net458),
    .A3(clknet_1_0__leaf_net465),
    .S0(net977),
    .S1(clknet_1_0__leaf_net473),
    .X(net474));
 sky130_fd_sc_hd__and3b_1 c592 (.A_N(clknet_1_1__leaf_net350),
    .B(clknet_1_0__leaf_net473),
    .C(clknet_1_1__leaf_net759),
    .X(net475));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net470),
    .A1(clknet_1_1__leaf_net465),
    .A2(net454),
    .A3(net231),
    .S0(clknet_1_0__leaf_net471),
    .S1(clknet_1_1__leaf_net759),
    .X(net476));
 sky130_fd_sc_hd__sdfbbp_1 c594 (.CLK(clknet_4_6_0_clk),
    .D(net4),
    .RESET_B(net462),
    .SCD(clknet_1_0__leaf_net261),
    .SCE(net928),
    .SET_B(net996),
    .Q(net478),
    .Q_N(net477));
 sky130_fd_sc_hd__or4_4 c595 (.A(net351),
    .B(clknet_1_0__leaf_net474),
    .C(net462),
    .D(clknet_1_1__leaf_net761),
    .X(net479));
 sky130_fd_sc_hd__mux4_4 c596 (.A0(clknet_1_0__leaf_net479),
    .A1(net956),
    .A2(net952),
    .A3(net928),
    .S0(net939),
    .S1(net748),
    .X(net480));
 sky130_fd_sc_hd__nor3b_1 c597 (.A(net858),
    .B(net250),
    .C_N(net477),
    .Y(net481));
 sky130_fd_sc_hd__nand3b_4 c598 (.A_N(net481),
    .B(clknet_1_0__leaf_net911),
    .C(net765),
    .Y(net482));
 sky130_fd_sc_hd__o2111ai_2 c599 (.A1(net819),
    .A2(net478),
    .B1(net942),
    .C1(net966),
    .D1(net765),
    .Y(net926));
 sky130_fd_sc_hd__a2111o_1 c600 (.A1(net970),
    .A2(net436),
    .B1(net890),
    .C1(net250),
    .D1(net747),
    .X(net483));
 sky130_fd_sc_hd__and4b_1 c601 (.A_N(net462),
    .B(net2),
    .C(net477),
    .D(net765),
    .X(net484));
 sky130_fd_sc_hd__o2111ai_1 c602 (.A1(clknet_1_1__leaf_net382),
    .A2(net477),
    .B1(net956),
    .C1(net883),
    .D1(net758),
    .Y(net485));
 sky130_fd_sc_hd__a2111oi_4 c603 (.A1(clknet_1_0__leaf_net482),
    .A2(net924),
    .B1(clknet_1_1__leaf_net382),
    .C1(clknet_1_1__leaf_net147),
    .D1(net765),
    .Y(net486));
 sky130_fd_sc_hd__o2111ai_2 c604 (.A1(net940),
    .A2(net478),
    .B1(net966),
    .C1(net924),
    .D1(net764),
    .Y(net487));
 sky130_fd_sc_hd__mux4_4 c605 (.A0(net437),
    .A1(clknet_1_1__leaf_net479),
    .A2(net481),
    .A3(net875),
    .S0(net758),
    .S1(net764),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net462),
    .A1(clknet_1_1__leaf_net474),
    .A2(net437),
    .A3(net928),
    .S0(net686),
    .S1(net764),
    .X(net489));
 sky130_fd_sc_hd__mux4_4 c607 (.A0(net359),
    .A1(clknet_1_0__leaf_net386),
    .A2(net747),
    .A3(clknet_1_1__leaf_net761),
    .S0(net766),
    .S1(net768),
    .X(net490));
 sky130_fd_sc_hd__sdfbbn_1 c608 (.CLK_N(clknet_4_6_0_clk),
    .D(net485),
    .RESET_B(clknet_1_0__leaf_net490),
    .SCD(net483),
    .SCE(net966),
    .SET_B(net103),
    .Q(net492),
    .Q_N(net491));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net437),
    .A1(net441),
    .A2(net491),
    .A3(net840),
    .S0(net4),
    .S1(net765),
    .X(net493));
 sky130_fd_sc_hd__a2111oi_4 c610 (.A1(net966),
    .A2(net940),
    .B1(clknet_1_1__leaf_net482),
    .C1(net686),
    .D1(net768),
    .Y(net494));
 sky130_fd_sc_hd__mux4_2 c611 (.A0(net492),
    .A1(clknet_1_1__leaf_net473),
    .A2(clknet_1_1__leaf_net474),
    .A3(net966),
    .S0(net929),
    .S1(clknet_1_1__leaf_net261),
    .X(net495));
 sky130_fd_sc_hd__a2111oi_4 c612 (.A1(net494),
    .A2(net484),
    .B1(clknet_1_1__leaf_net490),
    .C1(net957),
    .D1(net764),
    .Y(net496));
 sky130_fd_sc_hd__mux4_2 c613 (.A0(net478),
    .A1(net437),
    .A2(clknet_1_1__leaf_net496),
    .A3(clknet_1_1__leaf_net474),
    .S0(net491),
    .S1(clknet_1_0__leaf_net703),
    .X(net497));
 sky130_fd_sc_hd__sdfbbn_1 c614 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net474),
    .RESET_B(net483),
    .SCD(clknet_1_0__leaf_net381),
    .SCE(net942),
    .SET_B(clknet_1_1__leaf_net252),
    .Q(net499),
    .Q_N(net498));
 sky130_fd_sc_hd__mux4_2 c615 (.A0(clknet_1_0__leaf_net496),
    .A1(net492),
    .A2(clknet_1_1__leaf_net261),
    .A3(net498),
    .S0(net748),
    .S1(net749),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(clknet_1_1__leaf_net381),
    .A1(net929),
    .A2(net928),
    .A3(net233),
    .S0(net117),
    .S1(net754),
    .X(net501));
 sky130_fd_sc_hd__mux4_4 c617 (.A0(net250),
    .A1(net832),
    .A2(net949),
    .A3(net929),
    .S0(net883),
    .S1(net770),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net2),
    .A1(net878),
    .A2(net868),
    .A3(net952),
    .S0(net929),
    .S1(net771),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net834),
    .A1(net957),
    .A2(net843),
    .A3(net751),
    .S0(net752),
    .S1(net769),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c62 (.A0(net845),
    .A1(net3),
    .A2(net847),
    .A3(net849),
    .S0(net977),
    .S1(net976),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net928),
    .A1(net948),
    .A2(clknet_1_1__leaf_net386),
    .A3(net441),
    .S0(clknet_1_0__leaf_net880),
    .S1(net748),
    .X(net505));
 sky130_fd_sc_hd__mux4_4 c621 (.A0(clknet_1_1__leaf_net252),
    .A1(clknet_1_1__leaf_net147),
    .A2(net949),
    .A3(net105),
    .S0(net883),
    .S1(net751),
    .X(net506));
 sky130_fd_sc_hd__mux4_4 c622 (.A0(net32),
    .A1(clknet_1_1__leaf_net252),
    .A2(clknet_1_0__leaf_net880),
    .A3(net770),
    .S0(net771),
    .S1(net774),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net885),
    .A1(net928),
    .A2(net753),
    .A3(net872),
    .S0(net773),
    .S1(net1013),
    .X(net508));
 sky130_fd_sc_hd__mux4_4 c624 (.A0(net22),
    .A1(net288),
    .A2(net419),
    .A3(clknet_1_0__leaf_net409),
    .S0(net872),
    .S1(net772),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net871),
    .A1(net117),
    .A2(net877),
    .A3(net689),
    .S0(net751),
    .S1(net753),
    .X(net510));
 sky130_fd_sc_hd__mux4_4 c626 (.A0(clknet_1_0__leaf_net386),
    .A1(net510),
    .A2(net118),
    .A3(net924),
    .S0(net287),
    .S1(net882),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net5),
    .A1(net118),
    .A2(clknet_1_1__leaf_net409),
    .A3(net884),
    .S0(clknet_1_1__leaf_net911),
    .S1(net877),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net105),
    .A1(net360),
    .A2(net957),
    .A3(clknet_1_0__leaf_net511),
    .S0(net690),
    .S1(net769),
    .X(net876));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net246),
    .A1(net868),
    .A2(net878),
    .A3(net43),
    .S0(net873),
    .S1(net752),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c63 (.A0(net866),
    .A1(net849),
    .A2(net859),
    .A3(net858),
    .S0(net845),
    .S1(net977),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net475),
    .A1(net884),
    .A2(clknet_1_0__leaf_net876),
    .A3(net948),
    .S0(net754),
    .S1(net776),
    .X(net514));
 sky130_fd_sc_hd__mux4_2 c631 (.A0(net871),
    .A1(clknet_1_0__leaf_net386),
    .A2(clknet_1_0__leaf_net705),
    .A3(net771),
    .S0(net882),
    .S1(net773),
    .X(net515));
 sky130_fd_sc_hd__mux4_2 c632 (.A0(net419),
    .A1(clknet_1_1__leaf_net511),
    .A2(clknet_1_0__leaf_net386),
    .A3(net881),
    .S0(net710),
    .S1(net776),
    .X(net516));
 sky130_fd_sc_hd__mux4_4 c633 (.A0(net380),
    .A1(clknet_1_0__leaf_net409),
    .A2(clknet_1_0__leaf_net876),
    .A3(net957),
    .S0(clknet_1_0__leaf_net397),
    .S1(net771),
    .X(net517));
 sky130_fd_sc_hd__mux4_4 c634 (.A0(net32),
    .A1(clknet_1_1__leaf_net511),
    .A2(clknet_1_1__leaf_net705),
    .A3(net748),
    .S0(net776),
    .S1(net778),
    .X(net518));
 sky130_fd_sc_hd__mux4_4 c635 (.A0(clknet_1_0__leaf_net511),
    .A1(net22),
    .A2(net419),
    .A3(net767),
    .S0(net771),
    .S1(net778),
    .X(net519));
 sky130_fd_sc_hd__mux4_2 c636 (.A0(net233),
    .A1(net518),
    .A2(net957),
    .A3(net771),
    .S0(net778),
    .S1(clknet_1_0__leaf_net779),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net441),
    .A1(net520),
    .A2(net838),
    .A3(net754),
    .S0(net777),
    .S1(clknet_1_1__leaf_net779),
    .X(net521));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net853),
    .A1(net867),
    .A2(net864),
    .A3(net861),
    .S0(net849),
    .S1(net858),
    .X(net2));
 sky130_fd_sc_hd__or4_1 c65 (.A(net837),
    .B(net827),
    .C(net835),
    .D(net842),
    .X(net3));
 sky130_fd_sc_hd__or2_4 c66 (.A(net844),
    .B(net850),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 c660 (.A(net638),
    .X(net522));
 sky130_fd_sc_hd__inv_4 c661 (.A(net637),
    .Y(net523));
 sky130_fd_sc_hd__nand2_1 c662 (.A(net310),
    .B(net890),
    .Y(net524));
 sky130_fd_sc_hd__and2b_1 c663 (.A_N(net83),
    .B(net812),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_2 c664 (.A(net658),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_1 c665 (.A(net658),
    .X(net527));
 sky130_fd_sc_hd__inv_2 c666 (.A(net803),
    .Y(net528));
 sky130_fd_sc_hd__and2_1 c667 (.A(net812),
    .B(net964),
    .X(net529));
 sky130_fd_sc_hd__and2b_1 c668 (.A_N(net528),
    .B(net525),
    .X(net530));
 sky130_fd_sc_hd__or3_1 c669 (.A(net527),
    .B(net529),
    .C(net964),
    .X(net531));
 sky130_fd_sc_hd__or2_4 c67 (.A(net867),
    .B(net860),
    .X(net5));
 sky130_fd_sc_hd__or4_1 c670 (.A(net531),
    .B(net954),
    .C(net525),
    .D(net973),
    .X(net532));
 sky130_fd_sc_hd__inv_1 c671 (.A(net810),
    .Y(net533));
 sky130_fd_sc_hd__and4bb_1 c672 (.A_N(net532),
    .B_N(net420),
    .C(net523),
    .D(net964),
    .X(net534));
 sky130_fd_sc_hd__nand2b_2 c673 (.A_N(net531),
    .B(net964),
    .Y(net535));
 sky130_fd_sc_hd__or4b_1 c674 (.A(net529),
    .B(net531),
    .C(net535),
    .D_N(net965),
    .X(net536));
 sky130_fd_sc_hd__or2_1 c675 (.A(net528),
    .B(net530),
    .X(net537));
 sky130_fd_sc_hd__a2111oi_1 c676 (.A1(net523),
    .A2(net531),
    .B1(net537),
    .C1(net535),
    .D1(net964),
    .Y(net538));
 sky130_fd_sc_hd__nand2_1 c677 (.A(net530),
    .B(net529),
    .Y(net539));
 sky130_fd_sc_hd__and4b_1 c678 (.A_N(net539),
    .B(net964),
    .C(net535),
    .D(net536),
    .X(net540));
 sky130_fd_sc_hd__or3b_1 c679 (.A(net540),
    .B(net535),
    .C_N(net958),
    .X(net541));
 sky130_fd_sc_hd__or2_1 c68 (.A(net3),
    .B(net849),
    .X(net6));
 sky130_fd_sc_hd__o2111a_1 c680 (.A1(net967),
    .A2(net529),
    .B1(net208),
    .C1(net539),
    .D1(net964),
    .X(net542));
 sky130_fd_sc_hd__mux4_4 c681 (.A0(net536),
    .A1(net540),
    .A2(net529),
    .A3(net522),
    .S0(net307),
    .S1(net965),
    .X(net543));
 sky130_fd_sc_hd__nand2b_1 c682 (.A_N(net228),
    .B(net818),
    .Y(net544));
 sky130_fd_sc_hd__and3b_1 c683 (.A_N(net522),
    .B(net958),
    .C(net702),
    .X(net545));
 sky130_fd_sc_hd__or2_2 c684 (.A(clknet_1_1__leaf_net450),
    .B(net433),
    .X(net546));
 sky130_fd_sc_hd__nand3b_1 c685 (.A_N(net834),
    .B(clknet_1_0__leaf_net761),
    .C(clknet_1_0__leaf_net781),
    .Y(net547));
 sky130_fd_sc_hd__inv_1 c686 (.A(net804),
    .Y(net548));
 sky130_fd_sc_hd__nand3b_2 c687 (.A_N(net532),
    .B(net548),
    .C(net964),
    .Y(net549));
 sky130_fd_sc_hd__buf_4 c688 (.A(net810),
    .X(net550));
 sky130_fd_sc_hd__mux4_2 c689 (.A0(clknet_1_1__leaf_net453),
    .A1(net524),
    .A2(net549),
    .A3(net436),
    .S0(net834),
    .S1(net973),
    .X(net551));
 sky130_fd_sc_hd__and2_1 c69 (.A(net859),
    .B(net976),
    .X(net7));
 sky130_fd_sc_hd__nor3b_1 c690 (.A(net938),
    .B(clknet_1_0__leaf_net450),
    .C_N(net973),
    .Y(net552));
 sky130_fd_sc_hd__clkbuf_1 c691 (.A(net695),
    .X(net553));
 sky130_fd_sc_hd__inv_2 c692 (.A(net713),
    .Y(net554));
 sky130_fd_sc_hd__inv_2 c693 (.A(net695),
    .Y(net555));
 sky130_fd_sc_hd__inv_6 c694 (.A(net695),
    .Y(net556));
 sky130_fd_sc_hd__and3b_2 c695 (.A_N(net553),
    .B(net549),
    .C(clknet_1_1__leaf_net781),
    .X(net557));
 sky130_fd_sc_hd__nor3b_4 c696 (.A(net556),
    .B(net105),
    .C_N(clknet_1_0__leaf_net557),
    .Y(net558));
 sky130_fd_sc_hd__mux4_2 c697 (.A0(net548),
    .A1(clknet_1_0__leaf_net552),
    .A2(net556),
    .A3(clknet_1_0__leaf_net558),
    .S0(net549),
    .S1(net964),
    .X(net559));
 sky130_fd_sc_hd__or3b_1 c698 (.A(net541),
    .B(net958),
    .C_N(clknet_1_0__leaf_net558),
    .X(net560));
 sky130_fd_sc_hd__sdfbbp_1 c699 (.CLK(clknet_4_5_0_clk),
    .D(net546),
    .RESET_B(clknet_1_0__leaf_net560),
    .SCD(net228),
    .SCE(clknet_1_0__leaf_net551),
    .SET_B(net554),
    .Q(net562),
    .Q_N(net561));
 sky130_fd_sc_hd__and2_1 c70 (.A(net865),
    .B(net6),
    .X(net8));
 sky130_fd_sc_hd__mux4_2 c700 (.A0(net555),
    .A1(clknet_1_1__leaf_net560),
    .A2(net562),
    .A3(net550),
    .S0(net454),
    .S1(clknet_1_1__leaf_net557),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net549),
    .A1(clknet_1_0__leaf_net560),
    .A2(net561),
    .A3(clknet_1_0__leaf_net558),
    .S0(net545),
    .S1(net784),
    .X(net564));
 sky130_fd_sc_hd__mux4_4 c702 (.A0(net533),
    .A1(net562),
    .A2(net958),
    .A3(net549),
    .S0(clknet_1_0__leaf_net558),
    .S1(net785),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_2 c703 (.A(net695),
    .X(net566));
 sky130_fd_sc_hd__mux4_4 c704 (.A0(net958),
    .A1(net890),
    .A2(clknet_1_0__leaf_net467),
    .A3(clknet_1_0__leaf_net557),
    .S0(net968),
    .S1(net785),
    .X(net567));
 sky130_fd_sc_hd__a2111oi_2 c705 (.A1(net367),
    .A2(clknet_1_1__leaf_net558),
    .B1(net458),
    .C1(net566),
    .D1(net973),
    .Y(net568));
 sky130_fd_sc_hd__o2111a_4 c706 (.A1(clknet_1_1__leaf_net557),
    .A2(net362),
    .B1(clknet_1_0__leaf_net467),
    .C1(clknet_1_0__leaf_net473),
    .D1(net784),
    .X(net569));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net459),
    .RESET_B(clknet_1_0__leaf_net568),
    .SCD(clknet_1_0__leaf_net557),
    .SCE(net362),
    .SET_B(clknet_1_0__leaf_net569),
    .Q(net571),
    .Q_N(net570));
 sky130_fd_sc_hd__nor4b_1 c708 (.A(net537),
    .B(net842),
    .C(net965),
    .D_N(net958),
    .Y(net572));
 sky130_fd_sc_hd__mux4_2 c709 (.A0(net524),
    .A1(net469),
    .A2(clknet_1_0__leaf_net569),
    .A3(net360),
    .S0(net367),
    .S1(clknet_1_0__leaf_net467),
    .X(net573));
 sky130_fd_sc_hd__or2b_2 c71 (.A(net852),
    .B_N(net4),
    .X(net9));
 sky130_fd_sc_hd__and4b_1 c710 (.A_N(net362),
    .B(net458),
    .C(net87),
    .D(net965),
    .X(net574));
 sky130_fd_sc_hd__nor3_2 c711 (.A(net574),
    .B(net438),
    .C(clknet_1_1__leaf_net558),
    .Y(net575));
 sky130_fd_sc_hd__nand4_2 c712 (.A(clknet_1_1__leaf_net575),
    .B(clknet_1_1__leaf_net558),
    .C(net990),
    .D(net989),
    .Y(net576));
 sky130_fd_sc_hd__sedfxtp_2 c713 (.CLK(clknet_4_5_0_clk),
    .D(net231),
    .DE(clknet_1_0__leaf_net575),
    .SCD(clknet_1_0__leaf_net467),
    .SCE(net79),
    .Q(net577));
 sky130_fd_sc_hd__mux4_2 c714 (.A0(clknet_1_1__leaf_net558),
    .A1(clknet_1_1__leaf_net569),
    .A2(net566),
    .A3(clknet_1_0__leaf_net473),
    .S0(net87),
    .S1(net783),
    .X(net578));
 sky130_fd_sc_hd__sdfbbn_1 c715 (.CLK_N(clknet_4_5_0_clk),
    .D(net572),
    .RESET_B(clknet_1_0__leaf_net575),
    .SCD(net958),
    .SCE(clknet_1_1__leaf_net467),
    .SET_B(net784),
    .Q(net580),
    .Q_N(net579));
 sky130_fd_sc_hd__a2111o_1 c716 (.A1(net566),
    .A2(net571),
    .B1(clknet_1_0__leaf_net569),
    .C1(net965),
    .D1(net975),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(clknet_1_1__leaf_net581),
    .A1(net577),
    .A2(net580),
    .A3(net977),
    .S0(net535),
    .S1(clknet_1_0__leaf_net473),
    .X(net582));
 sky130_fd_sc_hd__mux4_4 c718 (.A0(net535),
    .A1(net567),
    .A2(net958),
    .A3(net458),
    .S0(net577),
    .S1(net965),
    .X(net583));
 sky130_fd_sc_hd__a2111o_4 c719 (.A1(net965),
    .A2(clknet_1_0__leaf_net581),
    .B1(net574),
    .C1(net783),
    .D1(net995),
    .X(net584));
 sky130_fd_sc_hd__or2_2 c72 (.A(net7),
    .B(net4),
    .X(net10));
 sky130_fd_sc_hd__sdfbbp_1 c720 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net583),
    .RESET_B(net1004),
    .SCD(net718),
    .SCE(net782),
    .SET_B(net995),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__clkinv_4 c455_7 (.A(clknet_1_1__leaf_net802),
    .Y(net984));
 sky130_fd_sc_hd__mux4_4 c722 (.A0(net468),
    .A1(net574),
    .A2(net585),
    .A3(net571),
    .S0(net709),
    .S1(net785),
    .X(net588));
 sky130_fd_sc_hd__mux4_4 c723 (.A0(net215),
    .A1(clknet_1_1__leaf_net557),
    .A2(net983),
    .A3(net959),
    .S0(clknet_1_0__leaf_net583),
    .S1(net570),
    .X(net589));
 sky130_fd_sc_hd__mux4_4 c724 (.A0(net577),
    .A1(net579),
    .A2(clknet_1_1__leaf_net583),
    .A3(net965),
    .S0(net982),
    .S1(net718),
    .X(net590));
 sky130_fd_sc_hd__mux4_4 c725 (.A0(net588),
    .A1(net578),
    .A2(clknet_1_1__leaf_net459),
    .A3(clknet_1_1__leaf_net569),
    .S0(clknet_1_0__leaf_net583),
    .S1(net788),
    .X(net591));
 sky130_fd_sc_hd__nand3_1 c726 (.A(net79),
    .B(net554),
    .C(net975),
    .Y(net592));
 sky130_fd_sc_hd__mux4_2 c727 (.A0(net436),
    .A1(net433),
    .A2(clknet_1_0__leaf_net583),
    .A3(clknet_1_1__leaf_net147),
    .S0(net585),
    .S1(net104),
    .X(net593));
 sky130_fd_sc_hd__a2111oi_4 c728 (.A1(net868),
    .A2(net968),
    .B1(net498),
    .C1(net832),
    .D1(net787),
    .Y(net594));
 sky130_fd_sc_hd__mux4_4 c729 (.A0(net977),
    .A1(clknet_1_1__leaf_net261),
    .A2(net965),
    .A3(net594),
    .S1(net788),
    .X(net595));
 sky130_fd_sc_hd__and2_1 c73 (.A(net6),
    .B(net8),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net868),
    .A1(net840),
    .A2(net550),
    .A3(net818),
    .S0(net855),
    .S1(net594),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net596),
    .A1(net554),
    .A2(net498),
    .A3(net594),
    .S0(net353),
    .S1(net999),
    .X(net597));
 sky130_fd_sc_hd__o2111ai_4 c732 (.A1(net592),
    .A2(net981),
    .B1(net436),
    .C1(clknet_1_1__leaf_net261),
    .D1(net554),
    .Y(net598));
 sky130_fd_sc_hd__a2111o_4 c733 (.A1(net499),
    .A2(net980),
    .B1(net526),
    .C1(net702),
    .D1(net763),
    .X(net599));
 sky130_fd_sc_hd__sdfbbn_1 c734 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net568),
    .RESET_B(net438),
    .SCD(net819),
    .SCE(net843),
    .SET_B(net999),
    .Q(net600));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net526),
    .A1(net586),
    .A2(net353),
    .A3(net499),
    .S0(net691),
    .S1(net975),
    .X(net601));
 sky130_fd_sc_hd__sdfbbn_1 c736 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net261),
    .RESET_B(net597),
    .SCD(net79),
    .SCE(net855),
    .SET_B(net1006),
    .Q(net603),
    .Q_N(net602));
 sky130_fd_sc_hd__nand4_1 c737 (.A(net580),
    .B(net603),
    .C(net594),
    .D(net788),
    .Y(net604));
 sky130_fd_sc_hd__a2111o_2 c738 (.A1(net600),
    .A2(net105),
    .B1(net603),
    .C1(net436),
    .D1(clknet_1_1__leaf_net467),
    .X(net605));
 sky130_fd_sc_hd__sdfbbp_1 c739 (.CLK(clknet_4_7_0_clk),
    .D(net594),
    .RESET_B(clknet_1_1__leaf_net467),
    .SCD(clknet_1_1__leaf_net261),
    .SCE(net603),
    .SET_B(net990),
    .Q(net606));
 sky130_fd_sc_hd__nand4_2 c74 (.A(net9),
    .B(net858),
    .C(net7),
    .D(net977),
    .Y(net12));
 sky130_fd_sc_hd__sdfbbn_2 c740 (.CLK_N(clknet_4_13_0_clk),
    .D(net487),
    .RESET_B(clknet_1_1__leaf_net147),
    .SCD(clknet_1_1__leaf_net467),
    .SCE(net889),
    .SET_B(net989),
    .Q(net608),
    .Q_N(net607));
 sky130_fd_sc_hd__sdfbbn_1 c741 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net583),
    .RESET_B(net601),
    .SCD(net499),
    .SCE(net550),
    .SET_B(net607),
    .Q(net609));
 sky130_fd_sc_hd__mux4_2 c742 (.A0(net606),
    .A1(net604),
    .A2(net840),
    .A3(net554),
    .S0(net979),
    .S1(net607),
    .X(net610));
 sky130_fd_sc_hd__a2111o_1 c743 (.A1(net610),
    .A2(net605),
    .B1(net609),
    .C1(net603),
    .D1(net978),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net499),
    .A1(net611),
    .A2(net608),
    .A3(clknet_1_1__leaf_net568),
    .S0(net602),
    .S1(clknet_1_0__leaf_net761),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net599),
    .A1(net487),
    .A2(net103),
    .A3(net607),
    .S0(net602),
    .S1(net790),
    .X(net613));
 sky130_fd_sc_hd__o2111a_1 c746 (.A1(net586),
    .A2(net608),
    .B1(net602),
    .C1(net554),
    .D1(net791),
    .X(net614));
 sky130_fd_sc_hd__nand4_4 c747 (.A(net359),
    .B(net614),
    .C(net608),
    .D(net762),
    .Y(net615));
 sky130_fd_sc_hd__mux4_4 c748 (.A0(net948),
    .A1(net968),
    .A2(net842),
    .A3(net615),
    .S0(net607),
    .S1(clknet_1_1__leaf_net780),
    .X(net616));
 sky130_fd_sc_hd__mux4_4 c749 (.A0(net360),
    .A1(net103),
    .A2(clknet_1_0__leaf_net397),
    .A3(clknet_1_1__leaf_net147),
    .S0(net550),
    .S1(clknet_1_0__leaf_net780),
    .X(net617));
 sky130_fd_sc_hd__nor2b_1 c75 (.A(net6),
    .B_N(net849),
    .Y(net13));
 sky130_fd_sc_hd__mux4_4 c750 (.A0(net608),
    .A1(net550),
    .A2(net832),
    .A3(clknet_1_1__leaf_net397),
    .S0(net615),
    .S1(net792),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net43),
    .A1(net513),
    .A2(net550),
    .A3(clknet_1_0__leaf_net618),
    .S0(net953),
    .S1(net792),
    .X(net619));
 sky130_fd_sc_hd__mux4_4 c752 (.A0(net957),
    .A1(clknet_1_1__leaf_net397),
    .A2(clknet_1_1__leaf_net616),
    .A3(net353),
    .S0(net615),
    .S1(net792),
    .X(net620));
 sky130_fd_sc_hd__mux4_2 c753 (.A0(net838),
    .A1(net615),
    .A2(clknet_1_1__leaf_net473),
    .A3(net225),
    .S0(net607),
    .S1(net792),
    .X(net621));
 sky130_fd_sc_hd__mux4_2 c754 (.A0(clknet_1_1__leaf_net618),
    .A1(clknet_1_1__leaf_net473),
    .A2(clknet_1_0__leaf_net397),
    .A3(net43),
    .S0(net615),
    .S1(clknet_1_0__leaf_net780),
    .X(net622));
 sky130_fd_sc_hd__mux4_2 c755 (.A0(clknet_1_1__leaf_net147),
    .A1(net554),
    .A2(net953),
    .A3(net615),
    .S0(net607),
    .S1(net792),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net619),
    .A1(net621),
    .A2(clknet_1_1__leaf_net397),
    .A3(clknet_1_1__leaf_net473),
    .S0(clknet_1_0__leaf_net616),
    .S1(net785),
    .X(net624));
 sky130_fd_sc_hd__mux4_2 c757 (.A0(net622),
    .A1(clknet_1_0__leaf_net616),
    .A2(net615),
    .A3(net788),
    .S0(net792),
    .S1(net794),
    .X(net625));
 sky130_fd_sc_hd__mux4_4 c758 (.A0(clknet_1_1__leaf_net625),
    .A1(net620),
    .A2(clknet_1_1__leaf_net397),
    .A3(net608),
    .S0(net792),
    .S1(net793),
    .X(net626));
 sky130_fd_sc_hd__mux4_2 c759 (.A0(net353),
    .A1(net842),
    .A2(net515),
    .A3(clknet_1_0__leaf_net626),
    .S0(net225),
    .S1(net794),
    .X(net627));
 sky130_fd_sc_hd__nand2b_1 c76 (.A_N(net827),
    .B(net10),
    .Y(net14));
 sky130_fd_sc_hd__mux4_2 c760 (.A0(net504),
    .A1(net627),
    .A2(clknet_1_0__leaf_net626),
    .A3(clknet_1_1__leaf_net703),
    .S0(net788),
    .S1(net793),
    .X(net628));
 sky130_fd_sc_hd__mux4_4 c761 (.A0(clknet_1_1__leaf_net628),
    .A1(clknet_1_1__leaf_net626),
    .A2(clknet_1_0__leaf_net625),
    .A3(net948),
    .S0(net792),
    .S1(net794),
    .X(net629));
 sky130_fd_sc_hd__mux4_2 c762 (.A0(net608),
    .A1(clknet_1_0__leaf_net628),
    .A2(clknet_1_1__leaf_net626),
    .A3(net615),
    .S0(net717),
    .S1(net788),
    .X(net630));
 sky130_fd_sc_hd__nor2_2 c77 (.A(net849),
    .B(net9),
    .Y(net15));
 sky130_fd_sc_hd__nor2b_1 c78 (.A(net856),
    .B_N(net7),
    .Y(net16));
 sky130_fd_sc_hd__and2b_2 c79 (.A_N(net822),
    .B(net7),
    .X(net17));
 sky130_fd_sc_hd__or2b_1 c80 (.A(net14),
    .B_N(net15),
    .X(net18));
 sky130_fd_sc_hd__nand2b_4 c81 (.A_N(net1),
    .B(net12),
    .Y(net19));
 sky130_fd_sc_hd__nor2_2 c82 (.A(net18),
    .B(net19),
    .Y(net20));
 sky130_fd_sc_hd__a2111o_1 c83 (.A1(net20),
    .A2(net10),
    .B1(net19),
    .C1(net17),
    .D1(net16),
    .X(net21));
 sky130_fd_sc_hd__and3b_4 c84 (.A_N(net839),
    .B(net20),
    .C(net17),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c85 (.A0(net20),
    .A1(net17),
    .A2(net15),
    .A3(net19),
    .S0(net7),
    .S1(net22),
    .X(net23));
 sky130_fd_sc_hd__o2111ai_1 c86 (.A1(net21),
    .A2(net23),
    .B1(net20),
    .C1(net4),
    .D1(net835),
    .Y(net24));
 sky130_fd_sc_hd__nand4b_4 c87 (.A_N(net24),
    .B(net14),
    .C(net20),
    .D(net15),
    .Y(net25));
 sky130_fd_sc_hd__and3b_1 c88 (.A_N(net21),
    .B(net2),
    .C(net19),
    .X(net26));
 sky130_fd_sc_hd__or3_4 c89 (.A(net841),
    .B(net860),
    .C(net835),
    .X(net27));
 sky130_fd_sc_hd__or3b_1 c90 (.A(net833),
    .B(net846),
    .C_N(net860),
    .X(net28));
 sky130_fd_sc_hd__and2b_2 c91 (.A_N(net841),
    .B(net11),
    .X(net29));
 sky130_fd_sc_hd__nor2_4 c92 (.A(net15),
    .B(net976),
    .Y(net891));
 sky130_fd_sc_hd__nand2_1 c93 (.A(net26),
    .B(net29),
    .Y(net30));
 sky130_fd_sc_hd__and2_4 c94 (.A(net860),
    .B(net891),
    .X(net31));
 sky130_fd_sc_hd__or2_2 c95 (.A(net9),
    .B(net30),
    .X(net32));
 sky130_fd_sc_hd__nand3b_1 c96 (.A_N(net27),
    .B(net21),
    .C(net32),
    .Y(net33));
 sky130_fd_sc_hd__or3_1 c97 (.A(net845),
    .B(net10),
    .C(net891),
    .X(net34));
 sky130_fd_sc_hd__and2_0 c98 (.A(net27),
    .B(net31),
    .X(net35));
 sky130_fd_sc_hd__nand2b_1 c99 (.A_N(net34),
    .B(net29),
    .Y(net36));
 sky130_fd_sc_hd__clkbuf_1 merge763 (.A(net693),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 merge764 (.A0(net12),
    .A1(net977),
    .A2(net124),
    .A3(net850),
    .S0(net96),
    .S1(clknet_1_1__leaf_net130),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 merge765 (.A0(net854),
    .A1(net124),
    .A2(net961),
    .A3(net38),
    .S0(net25),
    .S1(clknet_1_0__leaf_net147),
    .X(net633));
 sky130_fd_sc_hd__nor4b_2 merge766 (.A(net544),
    .B(clknet_1_1__leaf_net551),
    .C(net435),
    .D_N(net454),
    .Y(net634));
 sky130_fd_sc_hd__sdfbbp_1 merge767 (.CLK(clknet_4_4_0_clk),
    .D(net420),
    .SCD(net414),
    .SCE(net928),
    .SET_B(net413),
    .Q(net636),
    .Q_N(net421));
 sky130_fd_sc_hd__sdfrbp_1 merge768 (.CLK(clknet_4_4_0_clk),
    .D(net432),
    .RESET_B(net79),
    .SCD(net420),
    .SCE(net430),
    .Q(net638),
    .Q_N(net637));
 sky130_fd_sc_hd__sdfrbp_1 merge769 (.CLK(clknet_4_3_0_clk),
    .D(net251),
    .RESET_B(net352),
    .SCD(net111),
    .SCE(clknet_1_0__leaf_net252),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__or4_1 merge770 (.A(net71),
    .B(net208),
    .C(net308),
    .D(net193),
    .X(net641));
 sky130_fd_sc_hd__mux4_4 merge771 (.A0(net150),
    .A1(clknet_1_1__leaf_net252),
    .A2(net217),
    .A3(net259),
    .S0(net135),
    .S1(net929),
    .X(net642));
 sky130_fd_sc_hd__sdfbbn_1 merge772 (.CLK_N(clknet_4_6_0_clk),
    .D(net415),
    .RESET_B(net454),
    .SCD(net851),
    .SCE(net103),
    .SET_B(net942),
    .Q(net644),
    .Q_N(net643));
 sky130_fd_sc_hd__and4bb_1 merge773 (.A_N(net216),
    .B_N(net201),
    .C(net89),
    .D(net223),
    .X(net645));
 sky130_fd_sc_hd__mux4_2 merge774 (.A0(net238),
    .A1(net930),
    .A2(clknet_1_1__leaf_net252),
    .A3(net149),
    .S0(net136),
    .S1(net271),
    .X(net646));
 sky130_fd_sc_hd__mux4_4 merge775 (.A0(net55),
    .A1(net46),
    .A2(net62),
    .A3(net180),
    .S0(net178),
    .S1(net730),
    .X(net647));
 sky130_fd_sc_hd__mux4_4 merge776 (.A0(net94),
    .A1(net826),
    .A2(net830),
    .A3(net816),
    .S0(net95),
    .S1(net99),
    .X(net648));
 sky130_fd_sc_hd__mux4_4 merge777 (.A0(net236),
    .A1(net271),
    .A2(net918),
    .A3(net286),
    .S0(net5),
    .S1(net915),
    .X(net649));
 sky130_fd_sc_hd__o2111ai_1 merge778 (.A1(net223),
    .A2(net968),
    .B1(net811),
    .C1(net943),
    .D1(net201),
    .Y(net650));
 sky130_fd_sc_hd__and4bb_1 merge779 (.A_N(net337),
    .B_N(net230),
    .C(net220),
    .D(net103),
    .X(net651));
 sky130_fd_sc_hd__a2111o_2 merge780 (.A1(clknet_1_1__leaf_net552),
    .A2(net541),
    .B1(net547),
    .C1(net565),
    .D1(net784),
    .X(net652));
 sky130_fd_sc_hd__mux4_4 merge781 (.A0(net145),
    .A1(net142),
    .A2(clknet_1_0__leaf_net147),
    .A3(clknet_1_1__leaf_net245),
    .S0(net287),
    .S1(net271),
    .X(net653));
 sky130_fd_sc_hd__a2111o_1 merge782 (.A1(net60),
    .A2(net55),
    .B1(net139),
    .C1(net163),
    .D1(net42),
    .X(net654));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(net99),
    .A1(net1018),
    .A2(net98),
    .A3(net1012),
    .S0(net838),
    .S1(net201),
    .X(net655));
 sky130_fd_sc_hd__mux4_4 merge784 (.A0(net464),
    .A1(net103),
    .A2(net462),
    .A3(net127),
    .S0(net119),
    .S1(net975),
    .X(net656));
 sky130_fd_sc_hd__mux4_2 merge785 (.A0(net461),
    .A1(net928),
    .A2(net941),
    .A3(net573),
    .S0(clknet_1_0__leaf_net581),
    .S1(net718),
    .X(net657));
 sky130_fd_sc_hd__sdfrtn_1 merge786 (.CLK_N(clknet_4_4_0_clk),
    .D(net307),
    .RESET_B(net994),
    .SCD(net208),
    .SCE(net432),
    .Q(net658));
 sky130_fd_sc_hd__sdfbbn_1 merge787 (.CLK_N(clknet_4_8_0_clk),
    .D(clknet_1_1__leaf_net130),
    .RESET_B(net124),
    .SCD(net976),
    .SCE(net154),
    .SET_B(net41),
    .Q(net660),
    .Q_N(net659));
 sky130_fd_sc_hd__mux4_2 merge788 (.A0(net328),
    .A1(clknet_1_0__leaf_net350),
    .A2(clknet_1_0__leaf_net355),
    .A3(net260),
    .S0(net5),
    .S1(net132),
    .X(net661));
 sky130_fd_sc_hd__mux4_4 merge789 (.A0(net272),
    .A1(net271),
    .A2(net96),
    .A3(clknet_1_1__leaf_net130),
    .S0(net868),
    .S1(net739),
    .X(net662));
 sky130_fd_sc_hd__buf_6 merge790 (.A(net712),
    .X(net663));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net525),
    .A1(net958),
    .A2(net544),
    .A3(net430),
    .S0(net964),
    .S1(net527),
    .X(net664));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net869),
    .A1(net931),
    .A2(net854),
    .A3(net8),
    .S0(net139),
    .S1(clknet_1_0__leaf_net130),
    .X(net665));
 sky130_fd_sc_hd__mux4_2 merge793 (.A0(net214),
    .A1(net216),
    .A2(net220),
    .A3(net140),
    .S0(clknet_1_0__leaf_net261),
    .S1(net894),
    .X(net666));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net433),
    .A1(net424),
    .A2(net426),
    .A3(clknet_1_1__leaf_net322),
    .S0(net324),
    .S1(net326),
    .X(net667));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net179),
    .A1(net178),
    .A2(net169),
    .A3(clknet_1_1__leaf_net151),
    .S0(clknet_1_0__leaf_net147),
    .S1(net150),
    .X(net668));
 sky130_fd_sc_hd__mux4_4 merge796 (.A0(net97),
    .A1(net230),
    .A2(net224),
    .A3(net330),
    .S0(net220),
    .S1(net95),
    .X(net669));
 sky130_fd_sc_hd__mux4_4 merge797 (.A0(net1005),
    .A1(net256),
    .A2(clknet_1_0__leaf_net252),
    .A3(net198),
    .S0(net308),
    .S1(net205),
    .X(net670));
 sky130_fd_sc_hd__mux4_1 merge798 (.A0(net343),
    .A1(net959),
    .A2(clknet_1_0__leaf_net552),
    .A3(net219),
    .S0(net220),
    .S1(net1007),
    .X(net671));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net87),
    .A1(net531),
    .A2(net432),
    .A3(net545),
    .S0(net544),
    .S1(net958),
    .X(net672));
 sky130_fd_sc_hd__dfrbp_2 merge800 (.CLK(clknet_4_2_0_clk),
    .D(net648),
    .RESET_B(net655),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__dfrbp_1 merge801 (.CLK(clknet_4_11_0_clk),
    .D(net392),
    .RESET_B(net393),
    .Q(net675),
    .Q_N(net905));
 sky130_fd_sc_hd__dfrtn_1 merge802 (.CLK_N(clknet_4_11_0_clk),
    .D(net283),
    .RESET_B(net298),
    .Q(net915));
 sky130_fd_sc_hd__dfrtp_1 merge803 (.CLK(clknet_4_1_0_clk),
    .D(net323),
    .RESET_B(net641),
    .Q(net676));
 sky130_fd_sc_hd__dfrtp_1 merge804 (.CLK(clknet_4_6_0_clk),
    .D(net460),
    .RESET_B(net456),
    .Q(net677));
 sky130_fd_sc_hd__dfrtp_1 merge805 (.CLK(clknet_4_9_0_clk),
    .D(net375),
    .RESET_B(net378),
    .Q(net678));
 sky130_fd_sc_hd__nand2_2 merge806 (.A(net576),
    .B(net582),
    .Y(net679));
 sky130_fd_sc_hd__and2b_1 merge807 (.A_N(net185),
    .B(net186),
    .X(net680));
 sky130_fd_sc_hd__dfsbp_1 merge808 (.CLK(clknet_4_0_0_clk),
    .D(net209),
    .SET_B(net206),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__or2b_4 merge809 (.A(net131),
    .B_N(net128),
    .X(net683));
 sky130_fd_sc_hd__dfsbp_1 merge810 (.CLK(clknet_4_3_0_clk),
    .D(net340),
    .SET_B(net333),
    .Q(net685),
    .Q_N(net684));
 sky130_fd_sc_hd__dfstp_1 merge811 (.CLK(clknet_4_11_0_clk),
    .SET_B(net300),
    .Q(net301));
 sky130_fd_sc_hd__dfstp_1 merge812 (.CLK(clknet_4_13_0_clk),
    .D(net486),
    .SET_B(net493),
    .Q(net686));
 sky130_fd_sc_hd__dfstp_1 merge813 (.CLK(clknet_4_10_0_clk),
    .D(net927),
    .SET_B(net654),
    .Q(net902));
 sky130_fd_sc_hd__dlrbn_1 merge814 (.D(net167),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net173),
    .Q(net688),
    .Q_N(net687));
 sky130_fd_sc_hd__dlrbn_1 merge815 (.D(net507),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net509),
    .Q(net690),
    .Q_N(net689));
 sky130_fd_sc_hd__dlrbp_1 merge816 (.D(net593),
    .GATE(clknet_4_7_0_clk),
    .Q(net595),
    .Q_N(net691));
 sky130_fd_sc_hd__dlrbp_1 merge817 (.D(net452),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net667),
    .Q(net694),
    .Q_N(net693));
 sky130_fd_sc_hd__dlrtn_2 merge818 (.D(net634),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net652),
    .Q(net695));
 sky130_fd_sc_hd__dlrtn_1 merge819 (.D(net229),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net235),
    .Q(net696));
 sky130_fd_sc_hd__dlrtn_1 merge820 (.D(net412),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net425),
    .Q(net697));
 sky130_fd_sc_hd__dlrtp_1 merge821 (.D(net366),
    .GATE(clknet_4_6_0_clk),
    .Q(net368));
 sky130_fd_sc_hd__nor2_1 merge822 (.A(net630),
    .B(net623),
    .Y(net698));
 sky130_fd_sc_hd__dlrtp_2 merge823 (.D(net241),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net255),
    .Q(net923));
 sky130_fd_sc_hd__dlrtp_1 merge824 (.D(net270),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net266),
    .Q(net699));
 sky130_fd_sc_hd__edfxbp_1 merge825 (.CLK(clknet_4_8_0_clk),
    .D(net632),
    .DE(net653),
    .Q(net701),
    .Q_N(net700));
 sky130_fd_sc_hd__edfxtp_1 merge826 (.CLK(clknet_4_5_0_clk),
    .D(net534),
    .DE(net542),
    .Q(net702));
 sky130_fd_sc_hd__sdlclkp_1 merge827 (.CLK(clknet_4_13_0_clk),
    .GATE(net698),
    .SCE(net495),
    .GCLK(net703));
 sky130_fd_sc_hd__sdlclkp_2 merge828 (.CLK(clknet_4_14_0_clk),
    .GATE(net408),
    .SCE(net400),
    .GCLK(net704));
 sky130_fd_sc_hd__sdlclkp_4 merge829 (.CLK(clknet_4_15_0_clk),
    .GATE(net512),
    .SCE(net514),
    .GCLK(net705));
 sky130_fd_sc_hd__dfrbp_1 merge830 (.CLK(clknet_4_2_0_clk),
    .D(net645),
    .RESET_B(net683),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__or2b_1 merge831 (.A(net402),
    .B_N(net407),
    .X(net708));
 sky130_fd_sc_hd__dfrbp_1 merge832 (.CLK(clknet_4_6_0_clk),
    .D(net500),
    .RESET_B(net584),
    .Q(net710),
    .Q_N(net709));
 sky130_fd_sc_hd__dfrtn_1 merge833 (.CLK_N(clknet_4_9_0_clk),
    .D(net662),
    .RESET_B(net642),
    .Q(net711));
 sky130_fd_sc_hd__dfrtp_1 merge834 (.CLK(clknet_4_10_0_clk),
    .D(net190),
    .RESET_B(net680),
    .Q(net904));
 sky130_fd_sc_hd__dfrtp_4 merge835 (.CLK(clknet_4_0_0_clk),
    .D(net650),
    .RESET_B(net670),
    .Q(net712));
 sky130_fd_sc_hd__dfrtp_1 merge836 (.CLK(clknet_4_13_0_clk),
    .D(net598),
    .RESET_B(net405),
    .Q(net889));
 sky130_fd_sc_hd__dfsbp_2 merge837 (.CLK(clknet_4_3_0_clk),
    .D(net651),
    .SET_B(net671),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__dfsbp_1 merge838 (.CLK(clknet_4_8_0_clk),
    .D(net665),
    .SET_B(net174),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__dfstp_1 merge839 (.CLK(clknet_4_15_0_clk),
    .D(net629),
    .SET_B(net708),
    .Q(net717));
 sky130_fd_sc_hd__dfstp_1 merge840 (.CLK(clknet_4_7_0_clk),
    .D(net589),
    .SET_B(net679),
    .Q(net718));
 sky130_fd_sc_hd__dfxbp_1 s841 (.CLK(clknet_4_10_0_clk),
    .D(net63),
    .Q(net720),
    .Q_N(net719));
 sky130_fd_sc_hd__dfxbp_1 s842 (.CLK(clknet_4_10_0_clk),
    .D(net66),
    .Q(net896),
    .Q_N(net721));
 sky130_fd_sc_hd__dfxtp_1 s843 (.CLK(clknet_4_2_0_clk),
    .D(net108),
    .Q(net722));
 sky130_fd_sc_hd__dfxtp_1 s844 (.CLK(clknet_4_0_0_clk),
    .D(net109),
    .Q(net723));
 sky130_fd_sc_hd__dfxtp_1 s845 (.CLK(clknet_4_8_0_clk),
    .D(net123),
    .Q(net724));
 sky130_fd_sc_hd__dlclkp_1 s846 (.CLK(clknet_4_2_0_clk),
    .GATE(net126),
    .GCLK(net725));
 sky130_fd_sc_hd__dlclkp_2 s847 (.CLK(clknet_4_2_0_clk),
    .GATE(net129),
    .GCLK(net726));
 sky130_fd_sc_hd__dlclkp_4 s848 (.CLK(clknet_4_8_0_clk),
    .GATE(net146),
    .GCLK(net727));
 sky130_fd_sc_hd__dlxbn_1 s849 (.D(net155),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net729),
    .Q_N(net728));
 sky130_fd_sc_hd__dlxbn_1 s850 (.D(net156),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net731),
    .Q_N(net730));
 sky130_fd_sc_hd__dlxbp_1 s851 (.D(net172),
    .GATE(clknet_4_10_0_clk),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__dlxtn_1 s852 (.D(net210),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net734));
 sky130_fd_sc_hd__dlxtn_2 s853 (.D(net211),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net735));
 sky130_fd_sc_hd__dlxtn_4 s854 (.D(net232),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net894));
 sky130_fd_sc_hd__dlxtp_1 s855 (.D(net258),
    .GATE(clknet_4_9_0_clk),
    .Q(net887));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s856 (.D(net265),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net736));
 sky130_fd_sc_hd__dfxbp_1 s857 (.CLK(clknet_4_9_0_clk),
    .D(net269),
    .Q(net738),
    .Q_N(net737));
 sky130_fd_sc_hd__dfxbp_1 s858 (.CLK(clknet_4_9_0_clk),
    .D(net274),
    .Q(net740),
    .Q_N(net739));
 sky130_fd_sc_hd__dfxtp_1 s859 (.CLK(clknet_4_9_0_clk),
    .D(net277),
    .Q(net741));
 sky130_fd_sc_hd__dfxtp_1 s860 (.CLK(clknet_4_9_0_clk),
    .D(net278),
    .Q(net742));
 sky130_fd_sc_hd__dfxtp_1 s861 (.CLK(clknet_4_11_0_clk),
    .D(net290),
    .Q(net907));
 sky130_fd_sc_hd__dlclkp_1 s862 (.CLK(clknet_4_11_0_clk),
    .GATE(net299),
    .GCLK(net908));
 sky130_fd_sc_hd__dlclkp_2 s863 (.CLK(clknet_4_1_0_clk),
    .GATE(net315),
    .GCLK(net743));
 sky130_fd_sc_hd__dlclkp_4 s864 (.CLK(clknet_4_1_0_clk),
    .GATE(net320),
    .GCLK(net744));
 sky130_fd_sc_hd__dlxbn_1 s865 (.D(net321),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net746),
    .Q_N(net745));
 sky130_fd_sc_hd__dlxbn_2 s866 (.D(net347),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__dlxbp_1 s867 (.D(net369),
    .GATE(clknet_4_6_0_clk),
    .Q(net875),
    .Q_N(net749));
 sky130_fd_sc_hd__dlxtn_1 s868 (.D(net383),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net750));
 sky130_fd_sc_hd__dlxtn_2 s869 (.D(net389),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net883));
 sky130_fd_sc_hd__dlxtn_1 s870 (.D(net391),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net751));
 sky130_fd_sc_hd__dlxtp_1 s871 (.D(net394),
    .GATE(clknet_4_12_0_clk),
    .Q(net752));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s872 (.D(net395),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net753));
 sky130_fd_sc_hd__dfxbp_1 s873 (.CLK(clknet_4_14_0_clk),
    .D(net401),
    .Q(net872),
    .Q_N(net754));
 sky130_fd_sc_hd__dfxbp_1 s874 (.CLK(clknet_4_14_0_clk),
    .D(net404),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__dfxtp_1 s875 (.CLK(clknet_4_14_0_clk),
    .D(net406),
    .Q(net886));
 sky130_fd_sc_hd__dfxtp_1 s876 (.CLK(clknet_4_4_0_clk),
    .D(net429),
    .Q(net757));
 sky130_fd_sc_hd__dfxtp_2 s877 (.CLK(clknet_4_4_0_clk),
    .D(net431),
    .Q(net758));
 sky130_fd_sc_hd__dlclkp_1 s878 (.CLK(clknet_4_4_0_clk),
    .GATE(net444),
    .GCLK(net759));
 sky130_fd_sc_hd__dlclkp_2 s879 (.CLK(clknet_4_4_0_clk),
    .GATE(net451),
    .GCLK(net760));
 sky130_fd_sc_hd__dlclkp_4 s880 (.CLK(clknet_4_4_0_clk),
    .GATE(net455),
    .GCLK(net761));
 sky130_fd_sc_hd__dlxbn_1 s881 (.D(net476),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__dlxbn_2 s882 (.D(net480),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__dlxbp_1 s883 (.D(net488),
    .GATE(clknet_4_12_0_clk),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__dlxtn_1 s884 (.D(net489),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net768));
 sky130_fd_sc_hd__dlxtn_1 s885 (.D(net497),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net769));
 sky130_fd_sc_hd__dlxtn_1 s886 (.D(net501),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net770));
 sky130_fd_sc_hd__dlxtp_1 s887 (.D(net502),
    .GATE(clknet_4_12_0_clk),
    .Q(net771));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s888 (.D(net503),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net882));
 sky130_fd_sc_hd__dfxbp_1 s889 (.CLK(clknet_4_15_0_clk),
    .D(net505),
    .Q(net773),
    .Q_N(net772));
 sky130_fd_sc_hd__dfxbp_1 s890 (.CLK(clknet_4_14_0_clk),
    .D(net506),
    .Q(net775),
    .Q_N(net774));
 sky130_fd_sc_hd__dfxtp_1 s891 (.CLK(clknet_4_14_0_clk),
    .D(net508),
    .Q(net776));
 sky130_fd_sc_hd__dfxtp_1 s892 (.CLK(clknet_4_15_0_clk),
    .D(net516),
    .Q(net777));
 sky130_fd_sc_hd__dfxtp_1 s893 (.CLK(clknet_4_15_0_clk),
    .D(net517),
    .Q(net778));
 sky130_fd_sc_hd__dlclkp_1 s894 (.CLK(clknet_4_15_0_clk),
    .GATE(net519),
    .GCLK(net779));
 sky130_fd_sc_hd__dlclkp_2 s895 (.CLK(clknet_4_15_0_clk),
    .GATE(net521),
    .GCLK(net780));
 sky130_fd_sc_hd__dlclkp_4 s896 (.CLK(clknet_4_5_0_clk),
    .GATE(net543),
    .GCLK(net781));
 sky130_fd_sc_hd__dlxbn_1 s897 (.D(net559),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__dlxbn_2 s898 (.D(net563),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net785),
    .Q_N(net784));
 sky130_fd_sc_hd__dlxbp_1 s899 (.D(net564),
    .GATE(clknet_4_7_0_clk),
    .Q(net787),
    .Q_N(net786));
 sky130_fd_sc_hd__dlxtn_2 s900 (.D(net590),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net788));
 sky130_fd_sc_hd__dlxtn_1 s901 (.D(net591),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net789));
 sky130_fd_sc_hd__dlxtn_1 s902 (.D(net612),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net790));
 sky130_fd_sc_hd__dlxtp_1 s903 (.D(net613),
    .GATE(clknet_4_7_0_clk),
    .Q(net791));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s904 (.D(net617),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net792));
 sky130_fd_sc_hd__dfxbp_1 s905 (.CLK(clknet_4_13_0_clk),
    .D(net624),
    .Q(net794),
    .Q_N(net793));
 sky130_fd_sc_hd__dfxbp_1 s906 (.CLK(clknet_4_10_0_clk),
    .D(net633),
    .Q(net796),
    .Q_N(net795));
 sky130_fd_sc_hd__dfxtp_1 s907 (.CLK(clknet_4_9_0_clk),
    .D(net646),
    .Q(net797));
 sky130_fd_sc_hd__dfxtp_1 s908 (.CLK(clknet_4_10_0_clk),
    .D(net647),
    .Q(net798));
 sky130_fd_sc_hd__dfxtp_1 s909 (.CLK(clknet_4_11_0_clk),
    .D(net649),
    .Q(net799));
 sky130_fd_sc_hd__dlclkp_1 s910 (.CLK(clknet_4_3_0_clk),
    .GATE(net656),
    .GCLK(net800));
 sky130_fd_sc_hd__dlclkp_2 s911 (.CLK(clknet_4_7_0_clk),
    .GATE(net657),
    .GCLK(net801));
 sky130_fd_sc_hd__dlclkp_4 s912 (.CLK(clknet_4_9_0_clk),
    .GATE(net661),
    .GCLK(net802));
 sky130_fd_sc_hd__dlxbn_1 s913 (.D(net664),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net804),
    .Q_N(net803));
 sky130_fd_sc_hd__dlxbn_1 s914 (.D(net666),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net806),
    .Q_N(net805));
 sky130_fd_sc_hd__dlxbp_1 s915 (.D(net668),
    .GATE(clknet_4_11_0_clk),
    .Q(net808),
    .Q_N(net807));
 sky130_fd_sc_hd__dlxtn_2 s916 (.D(net669),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net809));
 sky130_fd_sc_hd__dlxtn_1 s917 (.D(net672),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net810));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net692));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net811));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net812));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net813));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(in13),
    .X(net814));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net816));
 sky130_fd_sc_hd__buf_2 input9 (.A(in16),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_8 input10 (.A(in17),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(in18),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in2),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(in21),
    .X(net823));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net824));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(in23),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(in24),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net827));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net828));
 sky130_fd_sc_hd__buf_1 input21 (.A(in27),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in28),
    .X(net830));
 sky130_fd_sc_hd__buf_1 input23 (.A(in29),
    .X(net831));
 sky130_fd_sc_hd__buf_4 input24 (.A(in3),
    .X(net832));
 sky130_fd_sc_hd__buf_1 input25 (.A(in30),
    .X(net833));
 sky130_fd_sc_hd__buf_4 input26 (.A(in31),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net835));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net837));
 sky130_fd_sc_hd__buf_4 input30 (.A(in35),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(in37),
    .X(net840));
 sky130_fd_sc_hd__buf_1 input33 (.A(in38),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_8 input34 (.A(in39),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(in4),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(in40),
    .X(net844));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net845));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net846));
 sky130_fd_sc_hd__buf_2 input39 (.A(in43),
    .X(net847));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net849));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net850));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(in48),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(in49),
    .X(net853));
 sky130_fd_sc_hd__buf_2 input46 (.A(in5),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(in50),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(in51),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(in52),
    .X(net857));
 sky130_fd_sc_hd__buf_4 input50 (.A(in53),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(in54),
    .X(net859));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net860));
 sky130_fd_sc_hd__buf_4 input53 (.A(in56),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in57),
    .X(net862));
 sky130_fd_sc_hd__buf_1 input55 (.A(in58),
    .X(net863));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net864));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(in6),
    .X(net865));
 sky130_fd_sc_hd__buf_1 input58 (.A(in60),
    .X(net866));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(in7),
    .X(net868));
 sky130_fd_sc_hd__buf_2 input61 (.A(in8),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in9),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net871),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net872),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net873),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net1025),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output67 (.A(net875),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(clknet_1_1__leaf_net876),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net877),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net878),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output71 (.A(net879),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(clknet_1_1__leaf_net880),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net881),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net882),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output75 (.A(net883),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net884),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net885),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net886),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net887),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net888),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output81 (.A(net889),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output82 (.A(net890),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net891),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net892),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(clknet_1_1__leaf_net893),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output86 (.A(net972),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net895),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net896),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net897),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net898),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net899),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net900),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(clknet_1_1__leaf_net901),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net902),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net903),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net904),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net905),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(clknet_1_1__leaf_net906),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net907),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(clknet_1_1__leaf_net908),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net909),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net910),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(clknet_1_1__leaf_net911),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output104 (.A(net932),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net913),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net933),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net915),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output108 (.A(net916),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net917),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net918),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net919),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net920),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net921),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net922),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output115 (.A(net923),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output116 (.A(net924),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net925),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output118 (.A(net926),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_1 wire119 (.A(net67),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net419),
    .X(net928));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(net244),
    .X(net929));
 sky130_fd_sc_hd__buf_1 wire122 (.A(net165),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_2 max_cap123 (.A(net932),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_2 max_cap124 (.A(net912),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_1 max_cap125 (.A(net914),
    .X(net933));
 sky130_fd_sc_hd__buf_1 wire126 (.A(net1022),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_1 max_cap127 (.A(net1023),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_2 max_cap128 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_2 wire129 (.A(net122),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_1 wire130 (.A(net538),
    .X(net938));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net314),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_2 max_cap132 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_2 wire133 (.A(net1021),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 fanout134 (.A(net246),
    .X(net942));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net199),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net313),
    .X(net944));
 sky130_fd_sc_hd__buf_1 max_cap137 (.A(net191),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_1 max_cap138 (.A(net44),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net50),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_2 max_cap140 (.A(net949),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_2 max_cap141 (.A(net42),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 max_cap142 (.A(net160),
    .X(net950));
 sky130_fd_sc_hd__buf_2 max_cap143 (.A(net342),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_2 max_cap144 (.A(net953),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_2 wire145 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_2 wire146 (.A(net955),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_2 max_cap147 (.A(net874),
    .X(net955));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net903),
    .X(net956));
 sky130_fd_sc_hd__buf_2 max_cap149 (.A(net469),
    .X(net957));
 sky130_fd_sc_hd__buf_2 fanout150 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net411),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(net962),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net113),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_2 max_cap155 (.A(net106),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net965),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net526),
    .X(net965));
 sky130_fd_sc_hd__buf_2 max_cap158 (.A(net481),
    .X(net966));
 sky130_fd_sc_hd__buf_1 max_cap159 (.A(net428),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_8 fanout160 (.A(net225),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net970),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net203),
    .X(net970));
 sky130_fd_sc_hd__buf_4 max_cap163 (.A(net752),
    .X(net971));
 sky130_fd_sc_hd__buf_12 fanout164 (.A(net894),
    .X(net972));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net734),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(net722),
    .X(net975));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(net863),
    .X(net976));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(net855),
    .X(net977));
 sky130_fd_sc_hd__inv_4 c721_1 (.A(clknet_1_1__leaf_net801),
    .Y(net978));
 sky130_fd_sc_hd__inv_4 net899_2 (.A(clknet_1_1__leaf_net801),
    .Y(net979));
 sky130_fd_sc_hd__inv_4 net899_3 (.A(clknet_1_1__leaf_net801),
    .Y(net980));
 sky130_fd_sc_hd__inv_4 net899_4 (.A(clknet_1_1__leaf_net801),
    .Y(net981));
 sky130_fd_sc_hd__inv_4 net899_5 (.A(clknet_1_0__leaf_net801),
    .Y(net982));
 sky130_fd_sc_hd__inv_4 net899_6 (.A(clknet_1_0__leaf_net801),
    .Y(net983));
 sky130_fd_sc_hd__clkinv_4 c455_8 (.A(clknet_1_0__leaf_net802),
    .Y(net985));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net802 (.A(net802),
    .X(clknet_0_net802));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net802 (.A(clknet_0_net802),
    .X(clknet_1_0__leaf_net802));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net802 (.A(clknet_0_net802),
    .X(clknet_1_1__leaf_net802));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net370 (.A(net370),
    .X(clknet_0_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_0__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net381 (.A(net381),
    .X(clknet_0_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_0__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_1__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net704 (.A(net704),
    .X(clknet_0_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net704 (.A(clknet_0_net704),
    .X(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net704 (.A(clknet_0_net704),
    .X(clknet_1_1__leaf_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net409 (.A(net409),
    .X(clknet_0_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_1__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net705 (.A(net705),
    .X(clknet_0_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_1__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net780 (.A(net780),
    .X(clknet_0_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net780 (.A(clknet_0_net780),
    .X(clknet_1_0__leaf_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net780 (.A(clknet_0_net780),
    .X(clknet_1_1__leaf_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net625 (.A(net625),
    .X(clknet_0_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net625 (.A(clknet_0_net625),
    .X(clknet_1_0__leaf_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net625 (.A(clknet_0_net625),
    .X(clknet_1_1__leaf_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net626 (.A(net626),
    .X(clknet_0_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net626 (.A(clknet_0_net626),
    .X(clknet_1_0__leaf_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net626 (.A(clknet_0_net626),
    .X(clknet_1_1__leaf_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net703 (.A(net703),
    .X(clknet_0_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net628 (.A(net628),
    .X(clknet_0_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net628 (.A(clknet_0_net628),
    .X(clknet_1_0__leaf_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net628 (.A(clknet_0_net628),
    .X(clknet_1_1__leaf_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net616 (.A(net616),
    .X(clknet_0_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_0__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_1__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net880 (.A(net880),
    .X(clknet_0_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net386 (.A(net386),
    .X(clknet_0_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net779 (.A(net779),
    .X(clknet_0_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net779 (.A(clknet_0_net779),
    .X(clknet_1_0__leaf_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net779 (.A(clknet_0_net779),
    .X(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net876 (.A(net876),
    .X(clknet_0_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net876 (.A(clknet_0_net876),
    .X(clknet_1_0__leaf_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net876 (.A(clknet_0_net876),
    .X(clknet_1_1__leaf_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net490 (.A(net490),
    .X(clknet_0_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net490 (.A(clknet_0_net490),
    .X(clknet_1_0__leaf_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net490 (.A(clknet_0_net490),
    .X(clknet_1_1__leaf_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net403 (.A(net403),
    .X(clknet_0_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_0__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_1__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net385 (.A(net385),
    .X(clknet_0_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_0__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_1__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net901 (.A(net901),
    .X(clknet_0_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net893 (.A(net893),
    .X(clknet_0_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net906 (.A(net906),
    .X(clknet_0_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net906 (.A(clknet_0_net906),
    .X(clknet_1_0__leaf_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net906 (.A(clknet_0_net906),
    .X(clknet_1_1__leaf_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net911 (.A(net911),
    .X(clknet_0_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net482 (.A(net482),
    .X(clknet_0_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_0__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_1__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net397 (.A(net397),
    .X(clknet_0_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_0__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_1__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net618 (.A(net618),
    .X(clknet_0_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net618 (.A(net986),
    .X(clknet_1_0__leaf_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net618 (.A(clknet_0_net618),
    .X(clknet_1_1__leaf_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net382 (.A(net382),
    .X(clknet_0_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_1__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net801 (.A(net801),
    .X(clknet_0_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net801 (.A(clknet_0_net801),
    .X(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net801 (.A(clknet_0_net801),
    .X(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net467 (.A(net467),
    .X(clknet_0_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_0__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net569 (.A(net569),
    .X(clknet_0_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net569 (.A(clknet_0_net569),
    .X(clknet_1_0__leaf_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net569 (.A(clknet_0_net569),
    .X(clknet_1_1__leaf_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net581 (.A(net581),
    .X(clknet_0_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_0__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_1__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net583 (.A(net583),
    .X(clknet_0_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_0__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_1__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net800 (.A(net800),
    .X(clknet_0_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_1__leaf_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net471 (.A(net471),
    .X(clknet_0_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_0__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_1__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net474 (.A(net474),
    .X(clknet_0_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_0__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_1__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net249 (.A(net249),
    .X(clknet_0_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_0__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_1__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net781 (.A(net781),
    .X(clknet_0_net781));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net781 (.A(clknet_0_net781),
    .X(clknet_1_0__leaf_net781));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net781 (.A(clknet_0_net781),
    .X(clknet_1_1__leaf_net781));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net557 (.A(net557),
    .X(clknet_0_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_0__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_1__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net558 (.A(net558),
    .X(clknet_0_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_0__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_1__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net575 (.A(net575),
    .X(clknet_0_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_1__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net568 (.A(net568),
    .X(clknet_0_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_0__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_1__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net560 (.A(net560),
    .X(clknet_0_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_0__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_1__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net761 (.A(net761),
    .X(clknet_0_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_0__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_1__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net760 (.A(net760),
    .X(clknet_0_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net760 (.A(clknet_0_net760),
    .X(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net760 (.A(clknet_0_net760),
    .X(clknet_1_1__leaf_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net759 (.A(net759),
    .X(clknet_0_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net453 (.A(net453),
    .X(clknet_0_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net453 (.A(clknet_0_net453),
    .X(clknet_1_0__leaf_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net453 (.A(clknet_0_net453),
    .X(clknet_1_1__leaf_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net551 (.A(net551),
    .X(clknet_0_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_0__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_1__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net450 (.A(net450),
    .X(clknet_0_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_0__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_1__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net552 (.A(net552),
    .X(clknet_0_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net552 (.A(clknet_0_net552),
    .X(clknet_1_0__leaf_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net552 (.A(clknet_0_net552),
    .X(clknet_1_1__leaf_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net744 (.A(net744),
    .X(clknet_0_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_1__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net371 (.A(net371),
    .X(clknet_0_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_0__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_1__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net322 (.A(net322),
    .X(clknet_0_net322));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net322 (.A(clknet_0_net322),
    .X(clknet_1_0__leaf_net322));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net322 (.A(clknet_0_net322),
    .X(clknet_1_1__leaf_net322));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net743 (.A(net743),
    .X(clknet_0_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net317 (.A(net317),
    .X(clknet_0_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_0__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_1__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net908 (.A(net908),
    .X(clknet_0_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_1__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net727 (.A(net727),
    .X(clknet_0_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net151 (.A(net151),
    .X(clknet_0_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net151 (.A(clknet_0_net151),
    .X(clknet_1_0__leaf_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net151 (.A(clknet_0_net151),
    .X(clknet_1_1__leaf_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net153 (.A(net153),
    .X(clknet_0_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net152 (.A(net152),
    .X(clknet_0_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net152 (.A(clknet_0_net152),
    .X(clknet_1_0__leaf_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net152 (.A(clknet_0_net152),
    .X(clknet_1_1__leaf_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net261 (.A(net261),
    .X(clknet_0_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net147 (.A(net147),
    .X(clknet_0_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net726 (.A(net726),
    .X(clknet_0_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_0__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_1__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net465 (.A(net465),
    .X(clknet_0_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_1__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net459 (.A(net459),
    .X(clknet_0_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_0__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_1__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net350 (.A(net350),
    .X(clknet_0_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_0__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_1__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net245 (.A(net245),
    .X(clknet_0_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net245 (.A(clknet_0_net245),
    .X(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net245 (.A(clknet_0_net245),
    .X(clknet_1_1__leaf_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net252 (.A(net252),
    .X(clknet_0_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net247 (.A(net247),
    .X(clknet_0_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net130 (.A(net130),
    .X(clknet_0_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_1__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net725 (.A(net725),
    .X(clknet_0_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_0__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_1__leaf_net725));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net1028),
    .X(net363));
 sky130_fd_sc_hd__or3_1 clone2 (.A(net974),
    .B(net969),
    .C(net988),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(clknet_0_net618),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_1 clone4 (.A(net894),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net332),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net787),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net702),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net253),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net724),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net735),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net967),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net786),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net758),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net875),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net736),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net789),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net207),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net733),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net231),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net681),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net677),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net254),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net785),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net676),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net848),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net732),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net696),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net447),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net219),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net775),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net740),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net135),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net678),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net904),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net100),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net796),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(net914),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(net314),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_1 max_cap3 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_1 wire4 (.A(net234),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_1 max_cap5 (.A(net44),
    .X(net1024));
 sky130_fd_sc_hd__buf_1 max_cap6 (.A(net874),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_1 fanout7 (.A(net969),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_1 fanout8 (.A(net974),
    .X(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_SCE (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SET_B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_SCE (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_C1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_Q_N (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_Q (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCD (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_Y (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_RESET_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_D (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_RESET_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_SCD (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_Q_N (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_Q (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_SCE (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_Q_N (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_Q (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_C1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_DE (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_D1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_Y (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_C (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_Y (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A_N (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net147_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_SCE (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_Y (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_X (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_SET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_SCE (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A3 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_SET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_Y (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_D (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_D (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_C (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_SET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A_N (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B_N (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_C1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_D1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_B_N (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_D (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_SCD (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Y (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_D (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_RESET_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_SCD (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A_N (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_B_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold19_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_D (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_SCE (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_C1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_Y (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B_N (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_X (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_C (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_C (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_D (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_D (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_Y (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_S0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_Y (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_C (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_SCD (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_C_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_C1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_C (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_Q (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net261_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_X (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_A_N (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_SET_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_D (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_D (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_D (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_SCD (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_X (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_Q_N (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_Q (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A_N (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_C_N (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Y (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_D (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_C1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A3 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Y (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_S1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_C (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_C (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_C (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_C1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A_N (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_D_N (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_SCD (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_C1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_X (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_C (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_X (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_C (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A_N (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCE (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_Q (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_C (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net397_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_X (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_C1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B_N (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_RESET_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_RESET_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_X (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_Y (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_Q_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_C (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_C_N (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_C1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_X (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_Y (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_RESET_B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_RESET_B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_DE (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_Y (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_SCD (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_RESET_B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_D_N (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_X (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_B_N (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B_N (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A2 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A_N (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_C (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_RESET_B (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_X (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_X (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_D1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_D (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_B1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_X (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_SCE (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_C1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_D1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_B (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_SET_B (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_Y (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A_N (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold7_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_Q (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_C1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_C (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_Q (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_Q (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_Q_N (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A_N (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_C (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_C (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_Y (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_s844_Q (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_C_N (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B_N (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_Q (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_Q (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_C1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_Q_N (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_Y (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_D (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_RESET_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_SCD (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCE (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_C (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A_N (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_Y (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A_N (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_C (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A_N (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_C (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_D1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A_N (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_C1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_SCE (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_SCD (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_Y (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A_N (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_C (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B_N (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A_N (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_SCD (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A_N (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_C1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A_N (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_C (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_C (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_D1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_C (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_SCE (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A_N (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_C (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_SCE (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_D1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_D (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_C (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_C (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_C1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_SCE (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_DE (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_SCD (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_C (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_D (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_C1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_SCE (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_SCE (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B_N (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_D (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_C (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_C1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_D1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_RESET_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A_N (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_C (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_C (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_C1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_C1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_Y (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_Q (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_RESET_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold14_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_Q (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_B_N (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_Q (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_C1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_Q (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_D (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_D (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_B1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_SCE (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_C (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_Y (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_C (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_C1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_C1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_Q (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_SCD (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_C (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_C (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_D (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_D (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_D1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_Y (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_Y (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_Q (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_C (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_SET_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_C1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCE (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_SCE (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_C (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_D (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_D (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap124_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap123_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_B1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_B1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B_N (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_SCE (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_SCE (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_SET_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_C_N (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_D_N (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_C (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_SET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_C1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_D1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_SCD (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap140_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap141_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap140_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap144_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire146_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire145_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap147_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire146_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap149_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_C1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCD (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_D_N (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_C_N (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_SCD (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_C_N (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A_N (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_D1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_C1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_D_N (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_B1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_C (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_C1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_D (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_D (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_C (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_C1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_D_N (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_C (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_C (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B_N (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_D1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_D1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_D1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_C_N (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_D (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_D_N (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SET_B (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_D1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_SCE (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_D (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_C1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_C (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_D1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_D1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_C_N (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_C (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_SCD (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_C1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_D (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s843_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s846_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_SLEEP_B (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s849_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s850_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net880_X (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net386_X (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCE (.DIODE(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_D1 (.DIODE(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_RESET_B (.DIODE(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_SCD (.DIODE(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net467_X (.DIODE(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B (.DIODE(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_C1 (.DIODE(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S1 (.DIODE(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net473_X (.DIODE(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(clknet_1_0__leaf_net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A2 (.DIODE(clknet_1_0__leaf_net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net552_X (.DIODE(clknet_1_0__leaf_net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_SCD (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCD (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net261_X (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_C1 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_D (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_SCD (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net261_X (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net147_A (.DIODE(clknet_0_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net147_A (.DIODE(clknet_0_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net147_X (.DIODE(clknet_0_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_S1 (.DIODE(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S0 (.DIODE(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net147_X (.DIODE(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_C1 (.DIODE(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_RESET_B (.DIODE(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net147_X (.DIODE(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_SCE (.DIODE(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_SCE (.DIODE(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCE (.DIODE(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A2 (.DIODE(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net252_X (.DIODE(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_SCD (.DIODE(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_SET_B (.DIODE(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A1 (.DIODE(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A2 (.DIODE(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net252_X (.DIODE(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_D_N (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_C (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_C (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_SCE (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_D1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_D1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SCE (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_D1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_D (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_C (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_D1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net103));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net335),
    .X(net1028));
 sky130_fd_sc_hd__or3_1 clone3 (.A(net1027),
    .B(net332),
    .C(net1026),
    .X(net1029));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
