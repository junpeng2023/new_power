module netlist_0 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input in52,
	input in53,
	input in54,
	input in55,
	input in56,
	input in57,
	input in58,
	input in59,
	input in60,
	input in61,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51,
	output out52,
	output out53,
	output out54,
	output out55,
	output out56,
	output out57,
	output out58,
	output out59,
	output out60,
	output out61
);


wire clk;
wire net893;
wire net892;
wire net890;
wire net889;
wire net885;
wire net882;
wire net881;
wire net880;
wire net878;
wire net877;
wire out20;
wire net887;
wire net875;
wire net871;
wire out17;
wire net866;
wire net865;
wire net864;
wire net863;
wire net862;
wire net860;
wire out3;
wire net857;
wire net854;
wire net853;
wire net851;
wire net850;
wire net849;
wire net848;
wire out38;
wire out29;
wire net846;
wire net844;
wire net842;
wire net841;
wire net837;
wire out0;
wire net834;
wire net833;
wire out54;
wire out4;
wire net832;
wire net831;
wire net829;
wire out31;
wire net827;
wire net835;
wire out11;
wire net825;
wire net843;
wire net823;
wire net822;
wire net821;
wire net820;
wire net819;
wire net818;
wire net817;
wire net816;
wire net815;
wire out8;
wire net814;
wire net813;
wire net812;
wire net811;
wire net810;
wire net807;
wire net805;
wire net804;
wire out15;
wire net802;
wire net801;
wire net800;
wire net795;
wire net793;
wire net792;
wire net791;
wire net789;
wire net787;
wire net786;
wire net785;
wire net784;
wire net808;
wire net781;
wire net780;
wire net777;
wire net869;
wire net776;
wire net775;
wire out12;
wire net774;
wire net773;
wire net772;
wire net771;
wire net770;
wire net769;
wire out49;
wire net766;
wire net765;
wire net764;
wire net763;
wire net762;
wire net759;
wire net755;
wire net754;
wire net753;
wire net752;
wire net751;
wire net750;
wire net748;
wire net790;
wire net747;
wire net745;
wire net744;
wire net743;
wire net741;
wire net740;
wire net739;
wire net738;
wire net735;
wire net732;
wire net731;
wire net730;
wire net729;
wire net728;
wire net726;
wire net725;
wire net724;
wire net722;
wire net720;
wire net719;
wire net717;
wire net716;
wire net715;
wire net714;
wire net712;
wire net711;
wire net708;
wire net706;
wire net705;
wire net704;
wire net703;
wire net701;
wire net699;
wire net692;
wire net690;
wire net895;
wire net299;
wire net688;
wire net686;
wire net684;
wire net683;
wire out57;
wire net503;
wire net679;
wire net671;
wire net669;
wire net668;
wire net370;
wire net667;
wire net664;
wire net694;
wire net659;
wire in6;
wire net656;
wire net652;
wire net622;
wire net651;
wire net304;
wire net645;
wire net641;
wire net637;
wire net632;
wire net665;
wire net631;
wire net629;
wire net74;
wire net628;
wire net3;
wire net627;
wire net447;
wire net626;
wire net624;
wire net506;
wire net623;
wire net620;
wire in49;
wire net619;
wire net879;
wire net798;
wire net46;
wire net615;
wire net347;
wire net100;
wire net288;
wire net614;
wire net165;
wire net613;
wire net20;
wire net612;
wire net638;
wire net428;
wire net610;
wire out25;
wire net608;
wire net1;
wire net424;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire net596;
wire net592;
wire net588;
wire net587;
wire in4;
wire net583;
wire net707;
wire net582;
wire net158;
wire net584;
wire net581;
wire net336;
wire net579;
wire net577;
wire net576;
wire net209;
wire net569;
wire in41;
wire net567;
wire net696;
wire net794;
wire in30;
wire net566;
wire net565;
wire net39;
wire net562;
wire net559;
wire net556;
wire net876;
wire net647;
wire net555;
wire net159;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire in55;
wire net550;
wire net867;
wire net710;
wire net544;
wire net539;
wire net534;
wire net532;
wire net271;
wire net530;
wire net617;
wire net306;
wire net537;
wire net369;
wire net528;
wire out13;
wire net525;
wire net523;
wire net872;
wire net520;
wire net519;
wire net516;
wire net672;
wire net514;
wire net78;
wire net508;
wire net721;
wire net504;
wire net224;
wire net573;
wire net499;
wire net674;
wire net496;
wire net495;
wire net494;
wire net888;
wire net179;
wire in39;
wire net453;
wire net493;
wire net788;
wire net472;
wire net492;
wire net897;
wire net479;
wire net491;
wire net295;
wire net490;
wire net489;
wire net856;
wire net487;
wire net486;
wire net478;
wire net474;
wire net473;
wire net468;
wire net540;
wire net202;
wire net465;
wire out7;
wire net462;
wire net469;
wire net471;
wire net461;
wire net546;
wire net749;
wire net460;
wire net454;
wire net44;
wire net117;
wire net689;
wire net859;
wire net858;
wire net648;
wire net452;
wire net449;
wire net448;
wire net498;
wire net700;
wire net446;
wire net680;
wire net88;
wire net691;
wire net444;
wire in59;
wire net110;
wire net442;
wire net441;
wire net609;
wire net440;
wire net128;
wire net439;
wire net147;
wire net438;
wire net797;
wire net433;
wire net432;
wire net419;
wire net431;
wire net430;
wire net618;
wire net429;
wire net427;
wire net809;
wire net426;
wire net673;
wire net425;
wire net423;
wire net183;
wire net531;
wire net421;
wire net52;
wire net170;
wire net420;
wire net450;
wire net418;
wire net415;
wire net414;
wire net276;
wire net413;
wire net330;
wire net252;
wire net412;
wire net411;
wire net826;
wire net517;
wire net677;
wire net410;
wire net409;
wire net685;
wire net407;
wire net662;
wire net405;
wire net836;
wire net607;
wire net526;
wire net404;
wire net29;
wire net403;
wire net383;
wire net663;
wire net402;
wire net106;
wire net572;
wire net401;
wire net847;
wire net399;
wire net398;
wire net476;
wire net855;
wire net396;
wire net172;
wire net395;
wire net779;
wire net698;
wire net839;
wire out23;
wire net391;
wire net693;
wire net884;
wire net443;
wire net557;
wire net345;
wire net527;
wire net488;
wire net390;
wire net646;
wire net389;
wire net513;
wire out14;
wire net501;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net184;
wire net131;
wire net380;
wire net379;
wire net260;
wire net616;
wire net378;
wire net543;
wire net38;
wire net377;
wire net376;
wire net625;
wire net373;
wire net598;
wire net374;
wire net676;
wire net861;
wire net372;
wire net371;
wire net368;
wire net475;
wire net408;
wire out26;
wire net367;
wire net366;
wire net365;
wire net364;
wire net782;
wire net601;
wire out35;
wire net363;
wire net360;
wire net660;
wire net838;
wire net359;
wire net397;
wire net357;
wire net356;
wire net510;
wire net355;
wire net570;
wire out2;
wire net521;
wire net353;
wire net590;
wire net507;
wire net351;
wire net746;
wire net350;
wire net547;
wire net511;
wire net451;
wire net13;
wire net343;
wire net89;
wire net666;
wire net340;
wire net339;
wire net337;
wire net406;
wire out19;
wire net458;
wire net538;
wire net244;
wire net334;
wire net333;
wire net332;
wire net331;
wire out43;
wire net328;
wire net327;
wire net119;
wire net325;
wire net324;
wire net321;
wire net535;
wire net320;
wire net542;
wire net139;
wire net318;
wire net316;
wire out9;
wire net335;
wire net315;
wire net313;
wire net505;
wire net199;
wire out27;
wire net294;
wire net319;
wire net312;
wire net309;
wire net417;
wire net302;
wire net298;
wire net286;
wire net153;
wire out61;
wire net296;
wire in24;
wire net358;
wire net127;
wire net697;
wire net293;
wire net305;
wire net594;
wire out39;
wire net292;
wire net500;
wire net445;
wire net230;
wire out22;
wire net303;
wire net291;
wire net201;
wire net422;
wire net289;
wire net595;
wire net384;
wire net482;
wire in25;
wire net272;
wire net142;
wire out10;
wire net589;
wire net278;
wire net761;
wire net274;
wire net643;
wire net273;
wire net114;
wire net270;
wire in17;
wire net267;
wire net644;
wire net266;
wire net459;
wire net463;
wire net0;
wire net297;
wire net280;
wire net102;
wire net799;
wire net151;
wire net275;
wire net264;
wire net657;
wire net591;
wire net196;
wire net262;
wire net217;
wire net261;
wire net21;
wire net257;
wire net62;
wire net109;
wire net254;
wire net203;
wire net253;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire in26;
wire net661;
wire net194;
wire net241;
wire net416;
wire net41;
wire net8;
wire net104;
wire out33;
wire in29;
wire net240;
wire net238;
wire net234;
wire out58;
wire net232;
wire net226;
wire out32;
wire net568;
wire net375;
wire net223;
wire net524;
wire net575;
wire net382;
wire net852;
wire net548;
wire net259;
wire net222;
wire net31;
wire net219;
wire net578;
wire net210;
wire net326;
wire net213;
wire net208;
wire out16;
wire net188;
wire net891;
wire net207;
wire net649;
wire net205;
wire net678;
wire net633;
wire net122;
wire net197;
wire net757;
wire in56;
wire net134;
wire out48;
wire net840;
wire net483;
wire net193;
wire net192;
wire net737;
wire net190;
wire net630;
wire in20;
wire net874;
wire net189;
wire net246;
wire net783;
wire net186;
wire net152;
wire net126;
wire net113;
wire net284;
wire net655;
wire net563;
wire net464;
wire net549;
wire net182;
wire net310;
wire net180;
wire out40;
wire net258;
wire net176;
wire net580;
wire net133;
wire net175;
wire net80;
wire net173;
wire in37;
wire net518;
wire net381;
wire net218;
wire net300;
wire net169;
wire net828;
wire net485;
wire net344;
wire net168;
wire net167;
wire net509;
wire net58;
wire net221;
wire net166;
wire net269;
wire net97;
wire net434;
wire net204;
wire net200;
wire net621;
wire net162;
wire out60;
wire net497;
wire out45;
wire net161;
wire net285;
wire net160;
wire net636;
wire net311;
wire net742;
wire net308;
wire out6;
wire out56;
wire net150;
wire in8;
wire net30;
wire out36;
wire net149;
wire net695;
wire net148;
wire net178;
wire net239;
wire net144;
wire net322;
wire net758;
wire net143;
wire out37;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net806;
wire net561;
wire net137;
wire net136;
wire net456;
wire net868;
wire net135;
wire net255;
wire net157;
wire net177;
wire net250;
wire net225;
wire net132;
wire net130;
wire in12;
wire net894;
wire net103;
wire net242;
wire net124;
wire out18;
wire net481;
wire net120;
wire net455;
wire net65;
wire net129;
wire net392;
wire net164;
wire net687;
wire net642;
wire net268;
wire in7;
wire net756;
wire net400;
wire net82;
wire net870;
wire net2;
wire net123;
wire net282;
wire net71;
wire net229;
wire in43;
wire net108;
wire net107;
wire net99;
wire net348;
wire net341;
wire in52;
wire net96;
wire net466;
wire net118;
wire net94;
wire net90;
wire net803;
wire net174;
wire net277;
wire net639;
wire net81;
wire in10;
wire net156;
wire net361;
wire net115;
wire net670;
wire in18;
wire net27;
wire net34;
wire net585;
wire net79;
wire net75;
wire net231;
wire net349;
wire net329;
wire net212;
wire net653;
wire in5;
wire net14;
wire net77;
wire net600;
wire net236;
wire net76;
wire in42;
wire net354;
wire in38;
wire net736;
wire net198;
wire net467;
wire net101;
wire net9;
wire net873;
wire net571;
wire net73;
wire net60;
wire net564;
wire net154;
wire net84;
wire net237;
wire net682;
wire in46;
wire net85;
wire net72;
wire net116;
wire net69;
wire net67;
wire in31;
wire net98;
wire net522;
wire net436;
wire net541;
wire net323;
wire net15;
wire net279;
wire net64;
wire net63;
wire net681;
wire net61;
wire net512;
wire net18;
wire out34;
wire net59;
wire net248;
wire net477;
wire net228;
wire net675;
wire net56;
wire out53;
wire net55;
wire net214;
wire net53;
wire in48;
wire net640;
wire net50;
wire net597;
wire out55;
wire net185;
wire net155;
wire net338;
wire net195;
wire out52;
wire net599;
wire net112;
wire net650;
wire net560;
wire net45;
wire net502;
wire net235;
wire net830;
wire net49;
wire in50;
wire net215;
wire net484;
wire net346;
wire net4;
wire net43;
wire net187;
wire in13;
wire net586;
wire net533;
wire net796;
wire net32;
wire net125;
wire net19;
wire in15;
wire net896;
wire net727;
wire net163;
wire in19;
wire net536;
wire net37;
wire net558;
wire in1;
wire net265;
wire out50;
wire net457;
wire net91;
wire net42;
wire net886;
wire net437;
wire in36;
wire out30;
wire net702;
wire net70;
wire net48;
wire net28;
wire net92;
wire net713;
wire net25;
wire in0;
wire net709;
wire net24;
wire out59;
wire out47;
wire net290;
wire net227;
wire net470;
wire in33;
wire net33;
wire net824;
wire net233;
wire net121;
wire net40;
wire in60;
wire net435;
wire net301;
wire net760;
wire net23;
wire net26;
wire net16;
wire net778;
wire net22;
wire net263;
wire net6;
wire net5;
wire net206;
wire in58;
wire net342;
wire net17;
wire in61;
wire net733;
wire net171;
wire in23;
wire in57;
wire net281;
wire net54;
wire in54;
wire in53;
wire net138;
wire net145;
wire net211;
wire out24;
wire in35;
wire in34;
wire net593;
wire in45;
wire net393;
wire net256;
wire net87;
wire net181;
wire net7;
wire out1;
wire net574;
wire net216;
wire in28;
wire in44;
wire net883;
wire in32;
wire net47;
wire net12;
wire in27;
wire in9;
wire net654;
wire net723;
wire net611;
wire net515;
wire net362;
wire in16;
wire net191;
wire out46;
wire net35;
wire net220;
wire in22;
wire net68;
wire in14;
wire net529;
wire in21;
wire net57;
wire net480;
wire net86;
wire net317;
wire in51;
wire net93;
wire in47;
wire in2;
wire net718;
wire net658;
wire net105;
wire in11;
wire net51;
wire net767;
wire net111;
wire net36;
wire net95;
wire net146;
wire net734;
wire net251;
wire net768;
wire net11;
wire net352;
wire net845;
wire net307;
wire net394;
wire net314;
wire in3;
sky130_fd_sc_hd__mux4_2 c62(
.A0(in51),
.A1(in57),
.A2(in46),
.A3(in44),
.S0(net3),
.S1(in48),
.X(net0)
);

sky130_fd_sc_hd__mux4_2 c63(
.A0(in52),
.A1(in45),
.A2(in54),
.A3(in49),
.S0(net3),
.S1(in46),
.X(net1)
);

sky130_fd_sc_hd__mux4_4 c64(
.A0(in58),
.A1(in56),
.A2(in61),
.A3(net3),
.S0(net0),
.S1(in46),
.X(net2)
);

sky130_fd_sc_hd__mux4_1 c65(
.A0(in36),
.A1(in23),
.A2(in28),
.A3(in21),
.S0(in10),
.S1(in22),
.X(net3)
);

sky130_fd_sc_hd__nand2_4 c66(
.A(in39),
.B(in32),
.Y(net4)
);

sky130_fd_sc_hd__nor3b_4 c67(
.A(in57),
.B(in48),
.C_N(net0),
.Y(net5)
);

sky130_fd_sc_hd__and2_2 c68(
.A(in35),
.B(in26),
.X(net6)
);

sky130_fd_sc_hd__buf_4 c69(
.A(net661),
.X(net7)
);

sky130_fd_sc_hd__clkinv_8 c70(
.A(net661),
.Y(net8)
);

sky130_fd_sc_hd__or2b_1 c71(
.A(net7),
.B_N(in10),
.X(net9)
);

sky130_fd_sc_hd__o211a_2 c72(
.A1(net8),
.A2(net5),
.B1(in58),
.C1(net1),
.X(net10)
);

sky130_fd_sc_hd__dlygate4sd3_1 c73(
.A(net669),
.X(net11)
);

sky130_fd_sc_hd__buf_16 c74(
.A(net769),
.X(net12)
);

sky130_fd_sc_hd__inv_12 c75(
.A(net788),
.Y(net13)
);

sky130_fd_sc_hd__o211a_4 c76(
.A1(net6),
.A2(net4),
.B1(net11),
.C1(net13),
.X(net14)
);

sky130_fd_sc_hd__mux4_1 c77(
.A0(net6),
.A1(in32),
.A2(in34),
.A3(net12),
.S0(net5),
.S1(net3),
.X(net15)
);

sky130_fd_sc_hd__o211a_2 c78(
.A1(net12),
.A2(net14),
.B1(in55),
.C1(in34),
.X(net16)
);

sky130_fd_sc_hd__clkinv_8 c79(
.A(net771),
.Y(net17)
);

sky130_fd_sc_hd__inv_8 c80(
.A(net669),
.Y(net18)
);

sky130_fd_sc_hd__and3b_1 c81(
.A_N(net9),
.B(net17),
.C(net740),
.X(net19)
);

sky130_fd_sc_hd__or2b_1 c82(
.A(in29),
.B_N(net740),
.X(net20)
);

sky130_fd_sc_hd__clkinv_4 c83(
.A(net790),
.Y(net21)
);

sky130_fd_sc_hd__or3_4 c84(
.A(net17),
.B(in21),
.C(net12),
.X(net22)
);

sky130_fd_sc_hd__inv_4 c85(
.A(net771),
.Y(net23)
);

sky130_fd_sc_hd__o211ai_4 c86(
.A1(net21),
.A2(net23),
.B1(net20),
.C1(net11),
.Y(net24)
);

sky130_fd_sc_hd__o211ai_4 c87(
.A1(net24),
.A2(net23),
.B1(net22),
.C1(net21),
.Y(net25)
);

sky130_fd_sc_hd__nand2_1 c88(
.A(net4),
.B(net14),
.Y(out30)
);

sky130_fd_sc_hd__inv_8 c89(
.A(net760),
.Y(net26)
);

sky130_fd_sc_hd__nor2_2 c90(
.A(net13),
.B(in53),
.Y(net27)
);

sky130_fd_sc_hd__dlygate4sd1_1 c91(
.A(net760),
.X(net28)
);

sky130_fd_sc_hd__nor2_4 c92(
.A(net17),
.B(net27),
.Y(net29)
);

sky130_fd_sc_hd__or3_2 c93(
.A(net7),
.B(net13),
.C(net29),
.X(net30)
);

sky130_fd_sc_hd__nand2b_2 c94(
.A_N(net27),
.B(in59),
.Y(net31)
);

sky130_fd_sc_hd__or2_1 c95(
.A(in52),
.B(in35),
.X(net32)
);

sky130_fd_sc_hd__clkbuf_2 c96(
.A(net805),
.X(net33)
);

sky130_fd_sc_hd__nor2_2 c97(
.A(net29),
.B(net26),
.Y(net34)
);

sky130_fd_sc_hd__nand2b_1 c98(
.A_N(net32),
.B(net33),
.Y(net35)
);

sky130_fd_sc_hd__or2b_2 c99(
.A(net33),
.B_N(in36),
.X(net36)
);

sky130_fd_sc_hd__nand2_2 c100(
.A(net20),
.B(net27),
.Y(net37)
);

sky130_fd_sc_hd__mux4_4 c101(
.A0(net35),
.A1(net36),
.A2(net37),
.A3(net28),
.S0(in35),
.S1(net33),
.X(net38)
);

sky130_fd_sc_hd__o211a_4 c102(
.A1(net37),
.A2(in36),
.B1(net33),
.C1(net35),
.X(net39)
);

sky130_fd_sc_hd__mux4_2 c103(
.A0(net26),
.A1(net36),
.A2(net33),
.A3(out30),
.S0(net39),
.S1(net34),
.X(net40)
);

sky130_fd_sc_hd__sdfrbp_1 c104(
.D(net39),
.RESET_B(net34),
.SCD(net33),
.SCE(net25),
.CLK(clk),
.Q(net42),
.Q_N(net41)
);

sky130_fd_sc_hd__inv_6 c105(
.A(net816),
.Y(net43)
);

sky130_fd_sc_hd__o211ai_2 c106(
.A1(in53),
.A2(net39),
.B1(net31),
.C1(net827),
.Y(net44)
);

sky130_fd_sc_hd__sdfrbp_2 c107(
.D(net31),
.RESET_B(net41),
.SCD(out30),
.SCE(net725),
.CLK(clk),
.Q(out47),
.Q_N(net45)
);

sky130_fd_sc_hd__mux4_2 c108(
.A0(net35),
.A1(net17),
.A2(net30),
.A3(net33),
.S0(net28),
.X(net46)
);

sky130_fd_sc_hd__sdfbbn_1 c109(
.D(net39),
.RESET_B(out47),
.SCD(net32),
.SCE(net41),
.SET_B(net725),
.CLK_N(clk),
.Q(net48),
.Q_N(net47)
);

sky130_fd_sc_hd__clkbuf_16 c110(
.A(net654),
.X(net49)
);

sky130_fd_sc_hd__nand2_2 c111(
.A(in29),
.B(net24),
.Y(net50)
);

sky130_fd_sc_hd__and3b_4 c112(
.A_N(net9),
.B(net11),
.C(net45),
.X(net51)
);

sky130_fd_sc_hd__and2b_1 c113(
.A_N(net43),
.B(in29),
.X(net52)
);

sky130_fd_sc_hd__or2_1 c114(
.A(in34),
.B(net45),
.X(net53)
);

sky130_fd_sc_hd__and2_1 c115(
.A(net24),
.B(net43),
.X(net54)
);

sky130_fd_sc_hd__nand2b_2 c116(
.A_N(net51),
.B(net52),
.Y(net55)
);

sky130_fd_sc_hd__nand2b_2 c117(
.A_N(in26),
.B(net43),
.Y(net56)
);

sky130_fd_sc_hd__o211a_4 c118(
.A1(net49),
.A2(net55),
.B1(net52),
.C1(out30),
.X(net57)
);

sky130_fd_sc_hd__sdfrtn_1 c119(
.D(net53),
.RESET_B(net48),
.SCD(in34),
.SCE(net55),
.CLK_N(clk),
.Q(net58)
);

sky130_fd_sc_hd__nor2b_1 c120(
.A(net32),
.B_N(net58),
.Y(net59)
);

sky130_fd_sc_hd__nor3_2 c121(
.A(net59),
.B(in32),
.C(net58),
.Y(net60)
);

sky130_fd_sc_hd__sdfrtp_1 c122(
.D(net52),
.RESET_B(net54),
.SCD(net60),
.SCE(net55),
.CLK(clk),
.Q(net61)
);

sky130_fd_sc_hd__inv_12 c123(
.A(net654),
.Y(out22)
);

sky130_fd_sc_hd__nand2_1 c124(
.A(net3),
.B(net51),
.Y(net62)
);

sky130_fd_sc_hd__o221ai_2 c125(
.A1(net62),
.A2(net59),
.B1(net58),
.B2(out30),
.C1(net61),
.Y(net63)
);

sky130_fd_sc_hd__mux4_2 c126(
.A0(net61),
.A1(in12),
.A2(in3),
.A3(net58),
.S0(in48),
.S1(net11),
.X(net64)
);

sky130_fd_sc_hd__o221a_1 c127(
.A1(net56),
.A2(net59),
.B1(net58),
.B2(in12),
.C1(net61),
.X(net65)
);

sky130_fd_sc_hd__mux4_1 c128(
.A0(net38),
.A1(net58),
.A2(net65),
.A3(net810),
.S0(net813),
.S1(net827),
.X(net66)
);

sky130_fd_sc_hd__clkinv_1 c129(
.A(net816),
.Y(net67)
);

sky130_fd_sc_hd__mux4_1 c130(
.A0(net50),
.A1(net67),
.A2(net62),
.A3(net65),
.S0(net51),
.S1(net58),
.X(net68)
);

sky130_fd_sc_hd__sdfbbn_2 c131(
.D(net62),
.RESET_B(net58),
.SCD(net54),
.SCE(net810),
.SET_B(net828),
.CLK_N(clk),
.Q(net70),
.Q_N(net69)
);

sky130_fd_sc_hd__and2_4 c132(
.A(in4),
.B(in7),
.X(net71)
);

sky130_fd_sc_hd__nand3b_2 c133(
.A_N(in17),
.B(in6),
.C(in15),
.Y(net72)
);

sky130_fd_sc_hd__nand2b_1 c134(
.A_N(net71),
.B(in17),
.Y(net73)
);

sky130_fd_sc_hd__o211ai_2 c135(
.A1(in4),
.A2(in18),
.B1(net71),
.C1(in3),
.Y(net74)
);

sky130_fd_sc_hd__or3_4 c136(
.A(in19),
.B(in8),
.C(net71),
.X(net75)
);

sky130_fd_sc_hd__or3b_2 c137(
.A(net75),
.B(in1),
.C_N(in12),
.X(net76)
);

sky130_fd_sc_hd__and2_2 c138(
.A(in13),
.B(in10),
.X(net77)
);

sky130_fd_sc_hd__inv_16 c139(
.A(net765),
.Y(net78)
);

sky130_fd_sc_hd__nor2_2 c140(
.A(in6),
.B(in2),
.Y(net79)
);

sky130_fd_sc_hd__o221ai_1 c141(
.A1(net75),
.A2(net73),
.B1(in18),
.B2(in7),
.C1(in9),
.Y(net80)
);

sky130_fd_sc_hd__or3_4 c142(
.A(in8),
.B(in16),
.C(net71),
.X(net81)
);

sky130_fd_sc_hd__inv_4 c143(
.A(net765),
.Y(net82)
);

sky130_fd_sc_hd__clkinv_1 c144(
.A(net749),
.Y(net83)
);

sky130_fd_sc_hd__mux4_1 c145(
.A0(in11),
.A1(net72),
.A2(net83),
.A3(net73),
.S0(net80),
.S1(in9),
.X(net84)
);

sky130_fd_sc_hd__or2_1 c146(
.A(net72),
.B(net763),
.X(net85)
);

sky130_fd_sc_hd__or2_1 c147(
.A(net82),
.B(in15),
.X(net86)
);

sky130_fd_sc_hd__or3_4 c148(
.A(net83),
.B(net85),
.C(net86),
.X(net87)
);

sky130_fd_sc_hd__clkinv_8 c149(
.A(net765),
.Y(net88)
);

sky130_fd_sc_hd__nand3b_2 c150(
.A_N(in15),
.B(net78),
.C(net83),
.Y(net89)
);

sky130_fd_sc_hd__nand3_1 c151(
.A(net74),
.B(net89),
.C(net86),
.Y(net90)
);

sky130_fd_sc_hd__o211a_1 c152(
.A1(net88),
.A2(net78),
.B1(net79),
.C1(net83),
.X(net91)
);

sky130_fd_sc_hd__sdfrtp_2 c153(
.D(net91),
.RESET_B(net90),
.SCD(net86),
.SCE(net81),
.CLK(clk),
.Q(net92)
);

sky130_fd_sc_hd__or2_4 c154(
.A(in43),
.B(in10),
.X(net93)
);

sky130_fd_sc_hd__or2_2 c155(
.A(in2),
.B(in23),
.X(net94)
);

sky130_fd_sc_hd__nor3b_2 c156(
.A(in30),
.B(net83),
.C_N(net94),
.Y(net95)
);

sky130_fd_sc_hd__nand3b_2 c157(
.A_N(in20),
.B(in30),
.C(net94),
.Y(net96)
);

sky130_fd_sc_hd__and2b_2 c158(
.A_N(net93),
.B(net94),
.X(net97)
);

sky130_fd_sc_hd__nor3_2 c159(
.A(net93),
.B(in40),
.C(net94),
.Y(net98)
);

sky130_fd_sc_hd__o211ai_1 c160(
.A1(net97),
.A2(net98),
.B1(in35),
.C1(net94),
.Y(net99)
);

sky130_fd_sc_hd__o211a_2 c161(
.A1(in18),
.A2(in42),
.B1(net98),
.C1(net94),
.X(net100)
);

sky130_fd_sc_hd__inv_12 c162(
.A(net759),
.Y(net101)
);

sky130_fd_sc_hd__mux4_2 c163(
.A0(in9),
.A1(in18),
.A2(net101),
.A3(net92),
.S0(net98),
.S1(net94),
.X(net102)
);

sky130_fd_sc_hd__o211a_1 c164(
.A1(net97),
.A2(in1),
.B1(net98),
.C1(net94),
.X(net103)
);

sky130_fd_sc_hd__o211ai_1 c165(
.A1(in25),
.A2(net103),
.B1(net99),
.C1(net94),
.Y(net104)
);

sky130_fd_sc_hd__buf_6 c166(
.A(net759),
.X(net105)
);

sky130_fd_sc_hd__clkbuf_2 c167(
.A(net771),
.X(net106)
);

sky130_fd_sc_hd__sdfbbp_1 c168(
.D(net105),
.RESET_B(net100),
.SCD(net101),
.SCE(net78),
.SET_B(net94),
.CLK(clk),
.Q(net108),
.Q_N(net107)
);

sky130_fd_sc_hd__nand3_4 c169(
.A(in33),
.B(net94),
.C(net765),
.Y(net109)
);

sky130_fd_sc_hd__o221a_2 c170(
.A1(net106),
.A2(net101),
.B1(net98),
.B2(net94),
.C1(net765),
.X(net110)
);

sky130_fd_sc_hd__o221a_1 c171(
.A1(net106),
.A2(net109),
.B1(net107),
.B2(net96),
.C1(net94),
.X(net111)
);

sky130_fd_sc_hd__sdfbbn_1 c172(
.D(net96),
.RESET_B(net105),
.SCD(net110),
.SCE(net109),
.SET_B(net94),
.CLK_N(clk),
.Q(net113),
.Q_N(net112)
);

sky130_fd_sc_hd__sdfbbn_2 c173(
.D(net110),
.RESET_B(net108),
.SCD(net113),
.SCE(net94),
.SET_B(net106),
.CLK_N(clk),
.Q(net115),
.Q_N(net114)
);

sky130_fd_sc_hd__mux4_1 c174(
.A0(net111),
.A1(net105),
.A2(net101),
.A3(net106),
.S0(net112),
.S1(net763),
.X(net116)
);

sky130_fd_sc_hd__mux4_2 c175(
.A0(net99),
.A1(net110),
.A2(in30),
.A3(net112),
.S0(net109),
.S1(net829),
.X(net117)
);

sky130_fd_sc_hd__clkinv_4 c176(
.A(net759),
.Y(net118)
);

sky130_fd_sc_hd__or2_1 c177(
.A(net108),
.B(net114),
.X(net119)
);

sky130_fd_sc_hd__nor2_2 c178(
.A(net119),
.B(net113),
.Y(net120)
);

sky130_fd_sc_hd__nor2b_1 c179(
.A(in49),
.B_N(net0),
.Y(net121)
);

sky130_fd_sc_hd__and2b_4 c180(
.A_N(in61),
.B(in58),
.X(net122)
);

sky130_fd_sc_hd__nand2b_2 c181(
.A_N(net83),
.B(net122),
.Y(net123)
);

sky130_fd_sc_hd__nor3_1 c182(
.A(in45),
.B(net123),
.C(net119),
.Y(net124)
);

sky130_fd_sc_hd__clkbuf_1 c183(
.A(net745),
.X(net125)
);

sky130_fd_sc_hd__or2_4 c184(
.A(net109),
.B(net125),
.X(out52)
);

sky130_fd_sc_hd__inv_1 c185(
.A(net820),
.Y(net126)
);

sky130_fd_sc_hd__buf_1 c186(
.A(net820),
.X(net127)
);

sky130_fd_sc_hd__dlygate4sd3_1 c187(
.A(net763),
.X(net128)
);

sky130_fd_sc_hd__nor2b_2 c188(
.A(net126),
.B_N(net123),
.Y(net129)
);

sky130_fd_sc_hd__mux4_4 c189(
.A0(net120),
.A1(net106),
.A2(in58),
.A3(net128),
.S0(net107),
.S1(net127),
.X(net130)
);

sky130_fd_sc_hd__and3b_2 c190(
.A_N(net128),
.B(net127),
.C(net94),
.X(net131)
);

sky130_fd_sc_hd__and2_1 c191(
.A(net131),
.B(net127),
.X(net132)
);

sky130_fd_sc_hd__inv_16 c192(
.A(net769),
.Y(net133)
);

sky130_fd_sc_hd__mux4_4 c193(
.A0(net125),
.A1(net77),
.A2(net124),
.A3(net132),
.S0(in23),
.S1(net112),
.X(net134)
);

sky130_fd_sc_hd__clkinv_4 c194(
.A(net763),
.Y(net135)
);

sky130_fd_sc_hd__or2_1 c195(
.A(net126),
.B(net830),
.X(net136)
);

sky130_fd_sc_hd__mux4_2 c196(
.A0(net133),
.A1(in50),
.A2(net136),
.A3(net83),
.S0(net98),
.S1(out52),
.X(net137)
);

sky130_fd_sc_hd__mux4_2 c197(
.A0(net132),
.A1(net122),
.A2(net136),
.A3(net127),
.S0(net135),
.S1(net830),
.X(net138)
);

sky130_fd_sc_hd__and3b_4 c198(
.A_N(net92),
.B(net115),
.C(net94),
.X(net139)
);

sky130_fd_sc_hd__o221ai_2 c199(
.A1(net139),
.A2(net22),
.B1(net71),
.B2(net136),
.C1(net96),
.Y(net140)
);

sky130_fd_sc_hd__buf_8 c200(
.A(net721),
.X(net141)
);

sky130_fd_sc_hd__clkbuf_16 c201(
.A(net810),
.X(net142)
);

sky130_fd_sc_hd__clkinv_8 c202(
.A(net789),
.Y(out46)
);

sky130_fd_sc_hd__and2_0 c203(
.A(net141),
.B(net740),
.X(net143)
);

sky130_fd_sc_hd__inv_1 c204(
.A(net790),
.Y(net144)
);

sky130_fd_sc_hd__and2b_4 c205(
.A_N(in27),
.B(net136),
.X(net145)
);

sky130_fd_sc_hd__nand3b_2 c206(
.A_N(net145),
.B(net127),
.C(net143),
.Y(net146)
);

sky130_fd_sc_hd__clkinv_4 c207(
.A(net777),
.Y(net147)
);

sky130_fd_sc_hd__nand3_4 c208(
.A(in55),
.B(net147),
.C(net830),
.Y(out55)
);

sky130_fd_sc_hd__clkbuf_1 c209(
.A(net721),
.X(net148)
);

sky130_fd_sc_hd__buf_1 c210(
.A(net743),
.X(net149)
);

sky130_fd_sc_hd__nand3b_2 c211(
.A_N(net136),
.B(net145),
.C(net148),
.Y(out36)
);

sky130_fd_sc_hd__sdfrtp_4 c212(
.D(net147),
.RESET_B(net141),
.SCD(net146),
.SCE(net5),
.CLK(clk),
.Q(net150)
);

sky130_fd_sc_hd__o211a_1 c213(
.A1(out55),
.A2(net115),
.B1(net144),
.C1(net830),
.X(net151)
);

sky130_fd_sc_hd__clkinv_2 c214(
.A(net771),
.Y(net152)
);

sky130_fd_sc_hd__inv_12 c215(
.A(net788),
.Y(net153)
);

sky130_fd_sc_hd__o211a_2 c216(
.A1(net148),
.A2(net150),
.B1(net149),
.C1(net151),
.X(out56)
);

sky130_fd_sc_hd__o211a_2 c217(
.A1(net150),
.A2(net146),
.B1(in28),
.C1(net153),
.X(net154)
);

sky130_fd_sc_hd__mux4_1 c218(
.A0(net152),
.A1(net149),
.A2(net146),
.A3(net141),
.S0(net153),
.S1(net721),
.X(net155)
);

sky130_fd_sc_hd__mux4_2 c219(
.A0(out36),
.A1(out56),
.A2(net136),
.A3(net146),
.S0(net721),
.S1(net832),
.X(net156)
);

sky130_fd_sc_hd__nand3_4 c220(
.A(in13),
.B(net127),
.C(net12),
.Y(net157)
);

sky130_fd_sc_hd__nor2b_2 c221(
.A(net29),
.B_N(in26),
.Y(out6)
);

sky130_fd_sc_hd__o211a_4 c222(
.A1(in12),
.A2(net28),
.B1(net157),
.C1(out36),
.X(net158)
);

sky130_fd_sc_hd__buf_2 c223(
.A(net813),
.X(net159)
);

sky130_fd_sc_hd__dlygate4sd1_1 c224(
.A(net804),
.X(net160)
);

sky130_fd_sc_hd__clkinv_2 c225(
.A(net760),
.Y(net161)
);

sky130_fd_sc_hd__or2b_2 c226(
.A(net12),
.B_N(net94),
.X(net162)
);

sky130_fd_sc_hd__sdfsbp_1 c227(
.D(net25),
.SCD(in34),
.SCE(net162),
.SET_B(net160),
.CLK(clk),
.Q(net164),
.Q_N(net163)
);

sky130_fd_sc_hd__o211ai_4 c228(
.A1(net30),
.A2(out55),
.B1(net25),
.C1(net14),
.Y(net165)
);

sky130_fd_sc_hd__o211ai_1 c229(
.A1(in26),
.A2(net29),
.B1(net163),
.C1(net2),
.Y(net166)
);

sky130_fd_sc_hd__o221ai_4 c230(
.A1(net143),
.A2(net19),
.B1(out47),
.B2(net160),
.C1(net28),
.Y(net167)
);

sky130_fd_sc_hd__o221ai_2 c231(
.A1(net28),
.A2(net160),
.B1(net47),
.B2(net12),
.C1(out55),
.Y(net168)
);

sky130_fd_sc_hd__nand2b_2 c232(
.A_N(net162),
.B(net769),
.Y(net169)
);

sky130_fd_sc_hd__sdfsbp_2 c233(
.D(out6),
.SCD(net127),
.SCE(net167),
.SET_B(net769),
.CLK(clk),
.Q(net171),
.Q_N(net170)
);

sky130_fd_sc_hd__buf_2 c234(
.A(net804),
.X(net172)
);

sky130_fd_sc_hd__sdfbbp_1 c235(
.D(in26),
.RESET_B(net157),
.SCD(out30),
.SCE(in54),
.SET_B(net729),
.CLK(clk),
.Q(net174),
.Q_N(net173)
);

sky130_fd_sc_hd__mux4_2 c236(
.A0(net157),
.A1(net22),
.A2(net171),
.A3(net162),
.S0(in48),
.S1(net172),
.X(net175)
);

sky130_fd_sc_hd__o221ai_2 c237(
.A1(in59),
.A2(net161),
.B1(net160),
.B2(net173),
.C1(net170),
.Y(net176)
);

sky130_fd_sc_hd__mux4_1 c238(
.A0(net23),
.A1(net174),
.A2(net167),
.A3(net160),
.S0(net169),
.S1(net176),
.X(net177)
);

sky130_fd_sc_hd__sdfstp_1 c239(
.D(net172),
.SCD(net164),
.SCE(net167),
.SET_B(net173),
.CLK(clk),
.Q(net178)
);

sky130_fd_sc_hd__nand2_1 c240(
.A(net174),
.B(net171),
.Y(net179)
);

sky130_fd_sc_hd__o221a_1 c241(
.A1(net179),
.A2(net178),
.B1(net159),
.B2(in48),
.C1(net779),
.X(out60)
);

sky130_fd_sc_hd__buf_1 c242(
.A(net798),
.X(net180)
);

sky130_fd_sc_hd__or3b_1 c243(
.A(net64),
.B(out47),
.C_N(out31),
.X(net181)
);

sky130_fd_sc_hd__and2_1 c244(
.A(net176),
.B(net168),
.X(net182)
);

sky130_fd_sc_hd__and3_4 c245(
.A(net14),
.B(net70),
.C(net64),
.X(net183)
);

sky130_fd_sc_hd__dlygate4sd1_1 c246(
.A(net798),
.X(out53)
);

sky130_fd_sc_hd__nor3b_2 c247(
.A(net160),
.B(net48),
.C_N(out53),
.Y(net184)
);

sky130_fd_sc_hd__clkinv_4 c248(
.A(net793),
.Y(net185)
);

sky130_fd_sc_hd__mux4_2 c249(
.A0(net164),
.A1(net54),
.A2(net180),
.A3(in21),
.S0(net160),
.S1(net14),
.X(net186)
);

sky130_fd_sc_hd__inv_12 c250(
.A(net789),
.Y(net187)
);

sky130_fd_sc_hd__mux4_4 c251(
.A0(net153),
.A1(net187),
.A2(net163),
.A3(net58),
.S0(net54),
.S1(net185),
.X(net188)
);

sky130_fd_sc_hd__o211a_1 c252(
.A1(net54),
.A2(net69),
.B1(net187),
.C1(out54),
.X(net189)
);

sky130_fd_sc_hd__and3b_2 c253(
.A_N(net187),
.B(net94),
.C(out54),
.X(net190)
);

sky130_fd_sc_hd__dfbbn_1 c254(
.D(net161),
.RESET_B(net185),
.SET_B(net183),
.CLK_N(clk),
.Q(net192),
.Q_N(net191)
);

sky130_fd_sc_hd__or3_1 c255(
.A(net14),
.B(out22),
.C(net787),
.X(out18)
);

sky130_fd_sc_hd__o221ai_2 c256(
.A1(net184),
.A2(net190),
.B1(net187),
.B2(out18),
.C1(out54),
.Y(net193)
);

sky130_fd_sc_hd__mux4_4 c257(
.A0(net190),
.A1(net64),
.A2(out18),
.A3(net47),
.S0(net183),
.S1(out54),
.X(net194)
);

sky130_fd_sc_hd__and3b_4 c258(
.A_N(net70),
.B(net77),
.C(net787),
.X(net195)
);

sky130_fd_sc_hd__buf_4 c259(
.A(net805),
.X(out48)
);

sky130_fd_sc_hd__mux4_2 c260(
.A0(net195),
.A1(net192),
.A2(out18),
.A3(net187),
.S0(net47),
.S1(net18),
.X(net196)
);

sky130_fd_sc_hd__mux4_2 c261(
.A0(in31),
.A1(net195),
.A2(out18),
.A3(net187),
.S0(net805),
.S1(out54),
.X(net197)
);

sky130_fd_sc_hd__mux4_2 c262(
.A0(net191),
.A1(net190),
.A2(out48),
.A3(net187),
.S0(out49),
.S1(net805),
.X(out40)
);

sky130_fd_sc_hd__o221a_4 c263(
.A1(net181),
.A2(net190),
.B1(net48),
.B2(out18),
.C1(out40),
.X(net198)
);

sky130_fd_sc_hd__nand2b_4 c264(
.A_N(in1),
.B(in7),
.Y(net199)
);

sky130_fd_sc_hd__and2_1 c265(
.A(in8),
.B(net85),
.X(net200)
);

sky130_fd_sc_hd__buf_12 c266(
.A(net735),
.X(net201)
);

sky130_fd_sc_hd__nand2b_4 c267(
.A_N(in15),
.B(net79),
.Y(net202)
);

sky130_fd_sc_hd__and2_0 c268(
.A(net202),
.B(net201),
.X(net203)
);

sky130_fd_sc_hd__buf_1 c269(
.A(net765),
.X(net204)
);

sky130_fd_sc_hd__inv_12 c270(
.A(net748),
.Y(net205)
);

sky130_fd_sc_hd__clkinv_4 c271(
.A(net735),
.Y(net206)
);

sky130_fd_sc_hd__inv_16 c272(
.A(net749),
.Y(net207)
);

sky130_fd_sc_hd__clkbuf_1 c273(
.A(net746),
.X(net208)
);

sky130_fd_sc_hd__or3b_2 c274(
.A(net202),
.B(net207),
.C_N(in5),
.X(net209)
);

sky130_fd_sc_hd__inv_16 c275(
.A(net751),
.Y(net210)
);

sky130_fd_sc_hd__nor3b_2 c276(
.A(net89),
.B(net208),
.C_N(net207),
.Y(net211)
);

sky130_fd_sc_hd__clkbuf_2 c277(
.A(net775),
.X(net212)
);

sky130_fd_sc_hd__inv_2 c278(
.A(net751),
.Y(net213)
);

sky130_fd_sc_hd__inv_6 c279(
.A(net734),
.Y(net214)
);

sky130_fd_sc_hd__and3_2 c280(
.A(net199),
.B(net207),
.C(net213),
.X(net215)
);

sky130_fd_sc_hd__mux4_1 c281(
.A0(net214),
.A1(net212),
.A2(net210),
.A3(in17),
.S0(net213),
.S1(net207),
.X(net216)
);

sky130_fd_sc_hd__sdfbbn_1 c282(
.D(net209),
.RESET_B(net216),
.SCD(net215),
.SCE(net213),
.SET_B(net212),
.CLK_N(clk),
.Q(net218),
.Q_N(net217)
);

sky130_fd_sc_hd__mux4_2 c283(
.A0(in14),
.A1(net213),
.A2(net215),
.A3(net217),
.S0(net200),
.S1(net209),
.X(net219)
);

sky130_fd_sc_hd__sdfbbn_2 c284(
.D(net202),
.RESET_B(net214),
.SCD(net217),
.SCE(net200),
.SET_B(net833),
.CLK_N(clk),
.Q(net221),
.Q_N(net220)
);

sky130_fd_sc_hd__mux4_1 c285(
.A0(net221),
.A1(net87),
.A2(net199),
.A3(net212),
.S0(net215),
.S1(net834),
.X(net222)
);

sky130_fd_sc_hd__nand2b_4 c286(
.A_N(net95),
.B(net215),
.Y(net223)
);

sky130_fd_sc_hd__nor2b_2 c287(
.A(in37),
.B_N(in23),
.Y(net224)
);

sky130_fd_sc_hd__mux4_1 c288(
.A0(net224),
.A1(net79),
.A2(net98),
.A3(net100),
.S0(net94),
.S1(net765),
.X(net225)
);

sky130_fd_sc_hd__dlygate4sd3_1 c289(
.A(net768),
.X(net226)
);

sky130_fd_sc_hd__or2b_4 c290(
.A(net79),
.B_N(net829),
.X(net227)
);

sky130_fd_sc_hd__nand2_4 c291(
.A(net93),
.B(net86),
.Y(net228)
);

sky130_fd_sc_hd__or2b_4 c292(
.A(net226),
.B_N(net224),
.X(net229)
);

sky130_fd_sc_hd__or3b_2 c293(
.A(in40),
.B(net212),
.C_N(net94),
.X(net230)
);

sky130_fd_sc_hd__and2b_1 c294(
.A_N(net101),
.B(in40),
.X(net231)
);

sky130_fd_sc_hd__nand2b_1 c295(
.A_N(net231),
.B(net212),
.Y(net232)
);

sky130_fd_sc_hd__or2b_1 c296(
.A(net231),
.B_N(net229),
.X(net233)
);

sky130_fd_sc_hd__o211ai_1 c297(
.A1(net232),
.A2(net230),
.B1(in24),
.C1(net94),
.Y(out58)
);

sky130_fd_sc_hd__o221a_1 c298(
.A1(net227),
.A2(in35),
.B1(net229),
.B2(net224),
.C1(net94),
.X(net234)
);

sky130_fd_sc_hd__clkinv_8 c299(
.A(net786),
.Y(net235)
);

sky130_fd_sc_hd__clkinv_4 c300(
.A(net768),
.Y(net236)
);

sky130_fd_sc_hd__o221a_1 c301(
.A1(net235),
.A2(net229),
.B1(net92),
.B2(net236),
.C1(net94),
.X(net237)
);

sky130_fd_sc_hd__buf_2 c302(
.A(net775),
.X(net238)
);

sky130_fd_sc_hd__clkbuf_4 c303(
.A(net734),
.X(net239)
);

sky130_fd_sc_hd__mux4_2 c304(
.A0(net100),
.A1(net236),
.A2(net233),
.A3(net217),
.S0(net231),
.S1(net224),
.X(net240)
);

sky130_fd_sc_hd__and2_1 c305(
.A(net218),
.B(net812),
.X(net241)
);

sky130_fd_sc_hd__or3b_4 c306(
.A(net241),
.B(net94),
.C_N(net812),
.X(net242)
);

sky130_fd_sc_hd__mux4_2 c307(
.A0(net242),
.A1(net237),
.A2(net238),
.A3(net235),
.S0(out58),
.S1(net224),
.X(net243)
);

sky130_fd_sc_hd__nand3_4 c308(
.A(in46),
.B(net224),
.C(net71),
.Y(net244)
);

sky130_fd_sc_hd__or3_4 c309(
.A(net235),
.B(net118),
.C(net831),
.X(net245)
);

sky130_fd_sc_hd__dlygate4sd1_1 c310(
.A(net768),
.X(net246)
);

sky130_fd_sc_hd__clkinv_8 c311(
.A(net748),
.Y(net247)
);

sky130_fd_sc_hd__buf_1 c312(
.A(net768),
.X(net248)
);

sky130_fd_sc_hd__mux4_4 c313(
.A0(net248),
.A1(net247),
.A2(net111),
.A3(net224),
.S0(out58),
.S1(net244),
.X(net249)
);

sky130_fd_sc_hd__mux4_4 c314(
.A0(net113),
.A1(net207),
.A2(net135),
.A3(net119),
.S0(net233),
.S1(in29),
.X(net250)
);

sky130_fd_sc_hd__o211a_1 c315(
.A1(net130),
.A2(in39),
.B1(net246),
.C1(net838),
.X(net251)
);

sky130_fd_sc_hd__or2_1 c316(
.A(net248),
.B(in48),
.X(net252)
);

sky130_fd_sc_hd__mux4_1 c317(
.A0(net233),
.A1(net224),
.A2(net215),
.A3(net113),
.S0(net831),
.S1(net838),
.X(net253)
);

sky130_fd_sc_hd__and2b_2 c318(
.A_N(net122),
.B(net819),
.X(net254)
);

sky130_fd_sc_hd__sdfstp_2 c319(
.D(net248),
.SCD(net244),
.SCE(net237),
.SET_B(net819),
.CLK(clk),
.Q(net255)
);

sky130_fd_sc_hd__nor3_4 c320(
.A(in31),
.B(in60),
.C(net831),
.Y(net256)
);

sky130_fd_sc_hd__nor3_4 c321(
.A(net118),
.B(net239),
.C(net838),
.Y(net257)
);

sky130_fd_sc_hd__nand3b_1 c322(
.A_N(net252),
.B(net255),
.C(net257),
.Y(net258)
);

sky130_fd_sc_hd__nor3_4 c323(
.A(net258),
.B(net255),
.C(net838),
.Y(out33)
);

sky130_fd_sc_hd__o211ai_2 c324(
.A1(net255),
.A2(net258),
.B1(in47),
.C1(net213),
.Y(net259)
);

sky130_fd_sc_hd__sdfstp_4 c325(
.D(net255),
.SCD(net237),
.SCE(net128),
.SET_B(net819),
.CLK(clk),
.Q(net260)
);

sky130_fd_sc_hd__sedfxbp_1 c326(
.D(net244),
.DE(net254),
.SCD(out33),
.SCE(net237),
.CLK(clk),
.Q(net262),
.Q_N(net261)
);

sky130_fd_sc_hd__sedfxbp_2 c327(
.D(net259),
.DE(net260),
.SCD(net256),
.SCE(net257),
.CLK(clk),
.Q(net264),
.Q_N(net263)
);

sky130_fd_sc_hd__and3b_4 c328(
.A_N(net260),
.B(net262),
.C(net119),
.X(net265)
);

sky130_fd_sc_hd__nor3b_2 c329(
.A(net206),
.B(net263),
.C_N(net831),
.Y(net266)
);

sky130_fd_sc_hd__nand3b_4 c330(
.A_N(net21),
.B(out46),
.C(net266),
.Y(net267)
);

sky130_fd_sc_hd__o211ai_4 c331(
.A1(net266),
.A2(out56),
.B1(net221),
.C1(net839),
.Y(net268)
);

sky130_fd_sc_hd__o221ai_4 c332(
.A1(in58),
.A2(net267),
.B1(net237),
.B2(net220),
.C1(net147),
.Y(net269)
);

sky130_fd_sc_hd__clkbuf_1 c333(
.A(net778),
.X(out32)
);

sky130_fd_sc_hd__o211a_4 c334(
.A1(net264),
.A2(net267),
.B1(net19),
.C1(net778),
.X(net270)
);

sky130_fd_sc_hd__buf_1 c335(
.A(net775),
.X(net271)
);

sky130_fd_sc_hd__o211a_2 c336(
.A1(in23),
.A2(net144),
.B1(net267),
.C1(net832),
.X(out34)
);

sky130_fd_sc_hd__clkinv_4 c337(
.A(net775),
.Y(net272)
);

sky130_fd_sc_hd__nand3_2 c338(
.A(net265),
.B(net267),
.C(net802),
.Y(net273)
);

sky130_fd_sc_hd__buf_12 c339(
.A(net786),
.X(net274)
);

sky130_fd_sc_hd__buf_12 c340(
.A(net778),
.X(net275)
);

sky130_fd_sc_hd__nand2_1 c341(
.A(net147),
.B(net275),
.Y(net276)
);

sky130_fd_sc_hd__nor3b_4 c342(
.A(net144),
.B(net115),
.C_N(net839),
.Y(net277)
);

sky130_fd_sc_hd__and2_1 c343(
.A(net276),
.B(net254),
.X(net278)
);

sky130_fd_sc_hd__o221a_2 c344(
.A1(net267),
.A2(net278),
.B1(net111),
.B2(in58),
.C1(out52),
.X(net279)
);

sky130_fd_sc_hd__clkbuf_8 c345(
.A(net776),
.X(net280)
);

sky130_fd_sc_hd__o221ai_1 c346(
.A1(net275),
.A2(net274),
.B1(net280),
.B2(net794),
.C1(net839),
.Y(net281)
);

sky130_fd_sc_hd__mux4_4 c347(
.A0(out58),
.A1(net275),
.A2(net281),
.A3(net19),
.S0(net280),
.S1(net802),
.X(net282)
);

sky130_fd_sc_hd__sdfbbp_1 c348(
.D(net221),
.RESET_B(net280),
.SCD(out52),
.SCE(net277),
.SET_B(net794),
.CLK(clk),
.Q(net284),
.Q_N(net283)
);

sky130_fd_sc_hd__mux4_1 c349(
.A0(net270),
.A1(net280),
.A2(net260),
.A3(out55),
.S0(net283),
.S1(net840),
.X(net285)
);

sky130_fd_sc_hd__mux4_4 c350(
.A0(net111),
.A1(net280),
.A2(net267),
.A3(out0),
.S0(net840),
.S1(net841),
.X(net286)
);

sky130_fd_sc_hd__mux4_2 c351(
.A0(net281),
.A1(net280),
.A2(net266),
.A3(net234),
.S0(net220),
.S1(net778),
.X(net287)
);

sky130_fd_sc_hd__clkinv_2 c352(
.A(net804),
.Y(out10)
);

sky130_fd_sc_hd__clkbuf_16 c353(
.A(net804),
.X(out39)
);

sky130_fd_sc_hd__and3_1 c354(
.A(net274),
.B(net141),
.C(net168),
.X(out1)
);

sky130_fd_sc_hd__mux4_2 c355(
.A0(net22),
.A1(net159),
.A2(out10),
.A3(net281),
.S0(out58),
.S1(net45),
.X(net288)
);

sky130_fd_sc_hd__clkbuf_1 c356(
.A(net808),
.X(out59)
);

sky130_fd_sc_hd__o221a_4 c357(
.A1(net141),
.A2(net175),
.B1(net38),
.B2(net94),
.C1(net842),
.X(net289)
);

sky130_fd_sc_hd__nand3b_1 c358(
.A_N(net213),
.B(net838),
.C(net842),
.Y(net290)
);

sky130_fd_sc_hd__o221ai_1 c359(
.A1(net290),
.A2(net18),
.B1(out32),
.B2(net729),
.C1(net842),
.Y(net291)
);

sky130_fd_sc_hd__sdfbbn_1 c360(
.D(net168),
.RESET_B(net291),
.SCD(out47),
.SCE(net159),
.SET_B(out58),
.CLK_N(clk),
.Q(net293),
.Q_N(net292)
);

sky130_fd_sc_hd__and3_4 c361(
.A(net19),
.B(out0),
.C(net842),
.X(net294)
);

sky130_fd_sc_hd__mux4_2 c362(
.A0(net293),
.A1(out60),
.A2(net178),
.A3(out46),
.S0(out56),
.S1(net835),
.X(net295)
);

sky130_fd_sc_hd__or3_2 c363(
.A(net271),
.B(in48),
.C(net42),
.X(net296)
);

sky130_fd_sc_hd__clkinv_2 c364(
.A(net760),
.Y(net297)
);

sky130_fd_sc_hd__nor3_1 c365(
.A(net19),
.B(net292),
.C(net290),
.Y(out61)
);

sky130_fd_sc_hd__and3b_2 c366(
.A_N(net290),
.B(net42),
.C(net94),
.X(net298)
);

sky130_fd_sc_hd__mux4_2 c367(
.A0(net273),
.A1(net18),
.A2(net169),
.A3(net291),
.S0(net774),
.S1(net844),
.X(net299)
);

sky130_fd_sc_hd__o221ai_1 c368(
.A1(net298),
.A2(net18),
.B1(net291),
.B2(out58),
.C1(out61),
.Y(net300)
);

sky130_fd_sc_hd__mux4_2 c369(
.A0(net18),
.A1(out58),
.A2(net290),
.A3(in48),
.S0(net19),
.S1(net845),
.X(net301)
);

sky130_fd_sc_hd__o221a_2 c370(
.A1(out52),
.A2(net291),
.B1(out34),
.B2(net774),
.C1(net812),
.X(net302)
);

sky130_fd_sc_hd__inv_4 c371(
.A(net813),
.Y(out37)
);

sky130_fd_sc_hd__mux4_1 c372(
.A0(net296),
.A1(net271),
.A2(net178),
.A3(net162),
.S0(out37),
.S1(net844),
.X(net303)
);

sky130_fd_sc_hd__mux4_1 c373(
.A0(out59),
.A1(out10),
.A2(net767),
.A3(net842),
.S0(net843),
.S1(net846),
.X(net304)
);

sky130_fd_sc_hd__mux4_4 c392(
.A0(net180),
.A1(out46),
.A2(in48),
.A3(net191),
.S0(out59),
.S1(net784),
.X(out45)
);

sky130_fd_sc_hd__mux4_1 c393(
.A0(net77),
.A1(net192),
.A2(out30),
.A3(out58),
.S0(out18),
.S1(out0),
.X(net305)
);

sky130_fd_sc_hd__mux4_4 c394(
.A0(net58),
.A1(in3),
.A2(net180),
.A3(out58),
.S0(net828),
.S1(out29),
.X(net306)
);

sky130_fd_sc_hd__mux4_1 c395(
.A0(net291),
.A1(net183),
.A2(out53),
.A3(out37),
.X(net307),
.S1(out29)
);

sky130_fd_sc_hd__nand2_1 c396(
.A(in7),
.B(net201),
.Y(net308)
);

sky130_fd_sc_hd__and2_1 c397(
.A(net201),
.B(net211),
.X(net309)
);

sky130_fd_sc_hd__inv_1 c398(
.A(net743),
.Y(net310)
);

sky130_fd_sc_hd__buf_16 c399(
.A(net719),
.X(net311)
);

sky130_fd_sc_hd__nand2_1 c400(
.A(net210),
.B(net199),
.Y(net312)
);

sky130_fd_sc_hd__inv_2 c401(
.A(net719),
.Y(net313)
);

sky130_fd_sc_hd__clkinv_4 c402(
.A(net732),
.Y(net314)
);

sky130_fd_sc_hd__or2b_4 c403(
.A(net211),
.B_N(net313),
.X(net315)
);

sky130_fd_sc_hd__inv_16 c404(
.A(net718),
.Y(net316)
);

sky130_fd_sc_hd__nor2_1 c405(
.A(net310),
.B(net218),
.Y(net317)
);

sky130_fd_sc_hd__sedfxtp_1 c406(
.D(net316),
.DE(net312),
.SCD(net313),
.SCE(net309),
.CLK(clk),
.Q(net318)
);

sky130_fd_sc_hd__sedfxtp_2 c407(
.D(net313),
.DE(net317),
.SCD(net315),
.SCE(net309),
.CLK(clk),
.Q(net319)
);

sky130_fd_sc_hd__mux4_1 c408(
.A0(net313),
.A1(net317),
.A2(net199),
.A3(net212),
.S0(net312),
.S1(net834),
.X(net320)
);

sky130_fd_sc_hd__or2b_4 c409(
.A(net312),
.B_N(net317),
.X(net321)
);

sky130_fd_sc_hd__inv_6 c410(
.A(net718),
.Y(net322)
);

sky130_fd_sc_hd__mux4_1 c411(
.A0(net216),
.A1(net321),
.A2(net311),
.A3(net314),
.S0(net319),
.S1(net309),
.X(net323)
);

sky130_fd_sc_hd__sedfxtp_4 c412(
.D(net311),
.DE(net322),
.SCD(net319),
.SCE(net309),
.CLK(clk),
.Q(net324)
);

sky130_fd_sc_hd__mux4_1 c413(
.A0(net321),
.A1(net313),
.A2(net316),
.A3(net320),
.S0(net317),
.S1(net319),
.X(net325)
);

sky130_fd_sc_hd__buf_6 c414(
.A(net746),
.X(net326)
);

sky130_fd_sc_hd__mux4_2 c415(
.A0(net314),
.A1(net321),
.A2(net310),
.A3(net200),
.S0(net319),
.S1(net309),
.X(net327)
);

sky130_fd_sc_hd__mux4_1 c416(
.A0(net326),
.A1(net324),
.A2(net309),
.A3(net818),
.S0(out38),
.S1(net847),
.X(net328)
);

sky130_fd_sc_hd__mux4_1 c417(
.A0(net322),
.A1(net311),
.A2(net71),
.A3(out38),
.S0(net847),
.S1(net848),
.X(net329)
);

sky130_fd_sc_hd__o211ai_2 c418(
.A1(net74),
.A2(net213),
.B1(net322),
.C1(net818),
.Y(net330)
);

sky130_fd_sc_hd__nor3_2 c419(
.A(net86),
.B(net236),
.C(net836),
.Y(out43)
);

sky130_fd_sc_hd__nor2b_2 c420(
.A(net226),
.B_N(net829),
.Y(net331)
);

sky130_fd_sc_hd__nor3_4 c421(
.A(net314),
.B(net331),
.C(net829),
.Y(net332)
);

sky130_fd_sc_hd__clkbuf_4 c422(
.A(net742),
.X(net333)
);

sky130_fd_sc_hd__and2b_4 c423(
.A_N(net314),
.B(net829),
.X(net334)
);

sky130_fd_sc_hd__o221a_4 c424(
.A1(in24),
.A2(net333),
.B1(net331),
.B2(net319),
.C1(net309),
.X(net335)
);

sky130_fd_sc_hd__nor2b_2 c425(
.A(net228),
.B_N(net322),
.Y(net336)
);

sky130_fd_sc_hd__nand2b_1 c426(
.A_N(net229),
.B(net236),
.Y(out19)
);

sky130_fd_sc_hd__buf_4 c427(
.A(net742),
.X(net337)
);

sky130_fd_sc_hd__o221ai_2 c428(
.A1(net236),
.A2(net326),
.B1(net310),
.B2(net739),
.C1(net847),
.Y(net338)
);

sky130_fd_sc_hd__mux4_1 c429(
.A0(net336),
.A1(out19),
.A2(net228),
.A3(net338),
.S0(net94),
.S1(net837),
.X(net339)
);

sky130_fd_sc_hd__mux4_1 c430(
.A0(net331),
.A1(net229),
.A2(net338),
.A3(out19),
.S0(out43),
.S1(net333),
.X(net340)
);

sky130_fd_sc_hd__nand3b_4 c431(
.A_N(in35),
.B(net338),
.C(net739),
.Y(net341)
);

sky130_fd_sc_hd__nor3b_1 c432(
.A(net341),
.B(net86),
.C_N(net849),
.Y(net342)
);

sky130_fd_sc_hd__mux4_1 c433(
.A0(net342),
.A1(in0),
.A2(net341),
.A3(net330),
.S0(net212),
.S1(in35),
.X(net343)
);

sky130_fd_sc_hd__mux4_2 c434(
.A0(net337),
.A1(net342),
.A2(out43),
.A3(net320),
.S0(net338),
.S1(net847),
.X(net344)
);

sky130_fd_sc_hd__mux4_4 c435(
.A0(out19),
.A1(net342),
.A2(net341),
.A3(net739),
.S0(net797),
.S1(net850),
.X(net345)
);

sky130_fd_sc_hd__mux4_4 c436(
.A0(in41),
.A1(net342),
.A2(net92),
.A3(net226),
.S0(net849),
.S1(net851),
.X(net346)
);

sky130_fd_sc_hd__mux4_4 c437(
.A0(net341),
.A1(net319),
.A2(net797),
.A3(net829),
.S0(net851),
.S1(net854),
.X(net347)
);

sky130_fd_sc_hd__mux4_1 c438(
.A0(net218),
.A1(net341),
.A2(net332),
.A3(net347),
.S0(net850),
.S1(net852),
.X(net348)
);

sky130_fd_sc_hd__mux4_2 c439(
.A0(net212),
.A1(net347),
.A2(net342),
.A3(net849),
.S0(net852),
.S1(net855),
.X(net349)
);

sky130_fd_sc_hd__or3b_4 c440(
.A(in22),
.B(net98),
.C_N(net254),
.X(net350)
);

sky130_fd_sc_hd__o221a_2 c441(
.A1(net247),
.A2(net207),
.B1(net333),
.B2(net739),
.C1(net850),
.X(net351)
);

sky130_fd_sc_hd__and3b_2 c442(
.A_N(net264),
.B(net245),
.C(net797),
.X(net352)
);

sky130_fd_sc_hd__sdfrbp_1 c443(
.D(in60),
.RESET_B(net215),
.SCD(net98),
.SCE(out33),
.CLK(clk),
.Q(out2),
.Q_N(net353)
);

sky130_fd_sc_hd__or3_1 c444(
.A(in39),
.B(net207),
.C(net334),
.X(net354)
);

sky130_fd_sc_hd__dlygate4sd1_1 c445(
.A(net784),
.X(net355)
);

sky130_fd_sc_hd__nand3b_2 c446(
.A_N(net355),
.B(net354),
.C(net850),
.Y(net356)
);

sky130_fd_sc_hd__o211ai_4 c447(
.A1(net351),
.A2(net98),
.B1(in0),
.C1(out2),
.Y(net357)
);

sky130_fd_sc_hd__nor3b_4 c448(
.A(net351),
.B(net835),
.C_N(net850),
.Y(net358)
);

sky130_fd_sc_hd__nand3_2 c449(
.A(net358),
.B(net354),
.C(net135),
.Y(net359)
);

sky130_fd_sc_hd__o211a_2 c450(
.A1(net359),
.A2(net215),
.B1(net355),
.C1(net263),
.X(net360)
);

sky130_fd_sc_hd__o221ai_4 c451(
.A1(net98),
.A2(net319),
.B1(net353),
.B2(net728),
.C1(net797),
.Y(net361)
);

sky130_fd_sc_hd__clkinv_16 c452(
.A(net784),
.Y(net362)
);

sky130_fd_sc_hd__sdfrbp_2 c453(
.D(in50),
.RESET_B(net320),
.SCD(out2),
.SCE(net361),
.CLK(clk),
.Q(out35),
.Q_N(net363)
);

sky130_fd_sc_hd__mux4_2 c454(
.A0(net256),
.A1(net119),
.A2(net362),
.A3(out35),
.S0(net353),
.S1(net856),
.X(net364)
);

sky130_fd_sc_hd__clkinv_8 c455(
.A(net776),
.Y(net365)
);

sky130_fd_sc_hd__buf_4 c456(
.A(net745),
.X(net366)
);

sky130_fd_sc_hd__o211ai_2 c457(
.A1(net326),
.A2(out2),
.B1(net94),
.C1(net728),
.Y(net367)
);

sky130_fd_sc_hd__mux4_1 c458(
.A0(net351),
.A1(net365),
.A2(in42),
.A3(net92),
.S0(net364),
.S1(net856),
.X(out26)
);

sky130_fd_sc_hd__mux4_4 c459(
.A0(net364),
.A1(net98),
.A2(in0),
.A3(net367),
.S0(net353),
.S1(out26),
.X(net368)
);

sky130_fd_sc_hd__mux4_1 c460(
.A0(net367),
.A1(net366),
.A2(net352),
.A3(in1),
.S0(out26),
.S1(net853),
.X(net369)
);

sky130_fd_sc_hd__mux4_1 c461(
.A0(net135),
.A1(net356),
.A2(net361),
.A3(net352),
.S0(net365),
.S1(out3),
.X(net370)
);

sky130_fd_sc_hd__nor3_1 c462(
.A(net365),
.B(net334),
.C(net832),
.Y(net371)
);

sky130_fd_sc_hd__nand3b_2 c463(
.A_N(in42),
.B(net371),
.C(net352),
.Y(net372)
);

sky130_fd_sc_hd__clkbuf_16 c464(
.A(net785),
.X(net373)
);

sky130_fd_sc_hd__and3b_2 c465(
.A_N(net371),
.B(net839),
.C(net854),
.X(net374)
);

sky130_fd_sc_hd__nor3_1 c466(
.A(net352),
.B(net284),
.C(in1),
.Y(net375)
);

sky130_fd_sc_hd__buf_2 c467(
.A(net785),
.X(net376)
);

sky130_fd_sc_hd__o211ai_2 c468(
.A1(net149),
.A2(in16),
.B1(in3),
.C1(in29),
.Y(net377)
);

sky130_fd_sc_hd__and3_1 c469(
.A(net377),
.B(net352),
.C(net812),
.X(net378)
);

sky130_fd_sc_hd__or3b_4 c470(
.A(net376),
.B(net8),
.C_N(net260),
.X(net379)
);

sky130_fd_sc_hd__clkinv_1 c471(
.A(net808),
.Y(net380)
);

sky130_fd_sc_hd__buf_4 c472(
.A(net800),
.X(net381)
);

sky130_fd_sc_hd__sdfbbn_2 c473(
.D(net373),
.RESET_B(net381),
.SCD(net5),
.SCE(net366),
.SET_B(net365),
.CLK_N(clk),
.Q(net383),
.Q_N(net382)
);

sky130_fd_sc_hd__o211a_4 c474(
.A1(net371),
.A2(net350),
.B1(net377),
.C1(net2),
.X(net384)
);

sky130_fd_sc_hd__inv_2 c475(
.A(net759),
.Y(net385)
);

sky130_fd_sc_hd__and3_4 c476(
.A(net385),
.B(net261),
.C(net818),
.X(net386)
);

sky130_fd_sc_hd__o221ai_4 c477(
.A1(net379),
.A2(net385),
.B1(net207),
.B2(net8),
.C1(net818),
.Y(net387)
);

sky130_fd_sc_hd__o221a_4 c478(
.A1(net272),
.A2(net387),
.B1(net381),
.B2(net385),
.C1(net841),
.X(net388)
);

sky130_fd_sc_hd__nor3_4 c479(
.A(net381),
.B(net246),
.C(net94),
.Y(out16)
);

sky130_fd_sc_hd__sdfbbp_1 c480(
.D(net388),
.RESET_B(net385),
.SCD(in0),
.SCE(net366),
.SET_B(net94),
.CLK(clk),
.Q(out7),
.Q_N(net389)
);

sky130_fd_sc_hd__o221a_1 c481(
.A1(net378),
.A2(net366),
.B1(net365),
.B2(net388),
.C1(net283),
.X(net390)
);

sky130_fd_sc_hd__mux4_2 c482(
.A0(net372),
.A1(net373),
.A2(net388),
.A3(net386),
.S0(net246),
.S1(net777),
.X(net391)
);

sky130_fd_sc_hd__mux4_2 c483(
.A0(net380),
.A1(net373),
.A2(out16),
.A3(net385),
.S0(net387),
.S1(net840),
.X(net392)
);

sky130_fd_sc_hd__o221a_2 c484(
.A1(net171),
.A2(net42),
.B1(net169),
.B2(net375),
.C1(net34),
.X(net393)
);

sky130_fd_sc_hd__o211a_2 c485(
.A1(net334),
.A2(out16),
.B1(net261),
.C1(net389),
.X(out23)
);

sky130_fd_sc_hd__o221a_4 c486(
.A1(out23),
.A2(net257),
.B1(in48),
.B2(net303),
.C1(net777),
.X(net394)
);

sky130_fd_sc_hd__sdfbbn_1 c487(
.D(out37),
.RESET_B(out1),
.SCD(net257),
.SCE(net71),
.SET_B(net812),
.CLK_N(clk),
.Q(net396),
.Q_N(net395)
);

sky130_fd_sc_hd__o221ai_4 c488(
.A1(net2),
.A2(net304),
.B1(net375),
.B2(net395),
.C1(net303),
.Y(net397)
);

sky130_fd_sc_hd__sdfrtn_1 c489(
.D(net375),
.RESET_B(net396),
.SCD(net34),
.SCE(net843),
.CLK_N(clk),
.Q(out27)
);

sky130_fd_sc_hd__mux4_4 c490(
.A0(net396),
.A1(out36),
.A2(out27),
.A3(net170),
.S0(net375),
.S1(net34),
.X(net398)
);

sky130_fd_sc_hd__o221a_1 c491(
.A1(net322),
.A2(out16),
.B1(out27),
.B2(in1),
.C1(net34),
.X(net399)
);

sky130_fd_sc_hd__o221a_4 c492(
.A1(net159),
.A2(net273),
.B1(net169),
.B2(net170),
.C1(net823),
.X(net400)
);

sky130_fd_sc_hd__sdfbbn_2 c493(
.D(net375),
.RESET_B(net372),
.SCD(net395),
.SCE(out33),
.SET_B(net823),
.CLK_N(clk),
.Q(out24),
.Q_N(net401)
);

sky130_fd_sc_hd__sdfbbp_1 c494(
.D(out39),
.RESET_B(net401),
.SCD(net392),
.SCE(out12),
.SET_B(net846),
.CLK(clk),
.Q(net403),
.Q_N(net402)
);

sky130_fd_sc_hd__mux4_2 c495(
.A0(net262),
.A1(net281),
.A2(in48),
.A3(in1),
.S0(net401),
.S1(net809),
.X(net404)
);

sky130_fd_sc_hd__mux4_4 c496(
.A0(net404),
.A1(out10),
.A2(out24),
.A3(net402),
.S0(net162),
.S1(out36),
.X(net405)
);

sky130_fd_sc_hd__mux4_4 c497(
.A0(net403),
.A1(net71),
.A2(out6),
.A3(net41),
.S0(net401),
.S1(out25),
.X(net406)
);

sky130_fd_sc_hd__mux4_4 c498(
.A0(net392),
.A1(net213),
.A2(net403),
.A3(net171),
.S0(net304),
.S1(out33),
.X(net407)
);

sky130_fd_sc_hd__mux4_2 c499(
.A0(net366),
.A1(out39),
.A2(net403),
.A3(out1),
.S0(net159),
.S1(net34),
.X(net408)
);

sky130_fd_sc_hd__mux4_4 c500(
.A0(net402),
.A1(in16),
.A2(net71),
.A3(out27),
.S0(net815),
.S1(net859),
.X(net409)
);

sky130_fd_sc_hd__sdfbbn_1 c501(
.D(net71),
.RESET_B(net2),
.SCD(out27),
.SCE(net159),
.SET_B(out24),
.CLK_N(clk),
.Q(net411),
.Q_N(net410)
);

sky130_fd_sc_hd__mux4_2 c502(
.A0(net304),
.A1(net410),
.A2(net366),
.A3(net303),
.S0(net784),
.S1(net859),
.X(net412)
);

sky130_fd_sc_hd__mux4_1 c503(
.A0(net411),
.A1(net409),
.A2(net401),
.A3(net809),
.S0(net859),
.S1(net860),
.X(net413)
);

sky130_fd_sc_hd__mux4_1 c504(
.A0(net413),
.A1(net411),
.A2(out27),
.A3(in48),
.S0(net859),
.S1(net860),
.X(net414)
);

sky130_fd_sc_hd__mux4_2 c505(
.A0(in1),
.A1(net409),
.A2(net404),
.A3(out24),
.S0(net375),
.S1(net410),
.X(net415)
);

sky130_fd_sc_hd__clkbuf_16 c528(
.A(net733),
.X(net416)
);

sky130_fd_sc_hd__and2_4 c529(
.A(net329),
.B(out38),
.X(net417)
);

sky130_fd_sc_hd__nor2_2 c530(
.A(net416),
.B(net848),
.Y(net418)
);

sky130_fd_sc_hd__clkinv_2 c531(
.A(net733),
.Y(net419)
);

sky130_fd_sc_hd__inv_16 c532(
.A(net776),
.Y(net420)
);

sky130_fd_sc_hd__and2_0 c533(
.A(in5),
.B(net420),
.X(net421)
);

sky130_fd_sc_hd__nand2b_1 c534(
.A_N(net420),
.B(net416),
.Y(net422)
);

sky130_fd_sc_hd__nor3_1 c535(
.A(net419),
.B(net319),
.C(net422),
.Y(net423)
);

sky130_fd_sc_hd__o211ai_4 c536(
.A1(net421),
.A2(net422),
.B1(net423),
.C1(in16),
.Y(net424)
);

sky130_fd_sc_hd__or2_2 c537(
.A(net420),
.B(net418),
.X(net425)
);

sky130_fd_sc_hd__and2_4 c538(
.A(net423),
.B(net421),
.X(net426)
);

sky130_fd_sc_hd__or2_2 c539(
.A(in16),
.B(net418),
.X(net427)
);

sky130_fd_sc_hd__buf_1 c540(
.A(net732),
.X(net428)
);

sky130_fd_sc_hd__and2_0 c541(
.A(net92),
.B(net418),
.X(net429)
);

sky130_fd_sc_hd__and2_0 c542(
.A(net428),
.B(net425),
.X(net430)
);

sky130_fd_sc_hd__buf_1 c543(
.A(net792),
.X(net431)
);

sky130_fd_sc_hd__nor3_2 c544(
.A(net431),
.B(net199),
.C(net418),
.Y(net432)
);

sky130_fd_sc_hd__inv_2 c545(
.A(net807),
.Y(net433)
);

sky130_fd_sc_hd__buf_2 c546(
.A(net806),
.X(net434)
);

sky130_fd_sc_hd__mux4_1 c547(
.A0(net434),
.A1(net422),
.A2(net419),
.A3(net421),
.S0(net424),
.S1(net429),
.X(net435)
);

sky130_fd_sc_hd__sdfbbn_2 c548(
.D(net425),
.RESET_B(net426),
.SCD(net308),
.SCE(net429),
.SET_B(net861),
.CLK_N(clk),
.Q(net437),
.Q_N(net436)
);

sky130_fd_sc_hd__nand3_1 c549(
.A(net432),
.B(net437),
.C(net861),
.Y(net438)
);

sky130_fd_sc_hd__or2_2 c550(
.A(net318),
.B(net847),
.X(net439)
);

sky130_fd_sc_hd__and2_1 c551(
.A(net436),
.B(net818),
.X(net440)
);

sky130_fd_sc_hd__inv_4 c552(
.A(net773),
.Y(net441)
);

sky130_fd_sc_hd__clkbuf_1 c553(
.A(net773),
.X(net442)
);

sky130_fd_sc_hd__nor2_1 c554(
.A(net439),
.B(net837),
.Y(net443)
);

sky130_fd_sc_hd__o221a_4 c555(
.A1(net441),
.A2(net310),
.B1(net94),
.B2(net427),
.C1(net436),
.X(net444)
);

sky130_fd_sc_hd__o211a_4 c556(
.A1(net440),
.A2(net427),
.B1(net338),
.C1(net836),
.X(net445)
);

sky130_fd_sc_hd__nor2_1 c557(
.A(net338),
.B(net440),
.Y(net446)
);

sky130_fd_sc_hd__sdfbbp_1 c558(
.D(net443),
.RESET_B(net338),
.SCD(net445),
.SCE(in31),
.SET_B(net849),
.CLK(clk),
.Q(net448),
.Q_N(net447)
);

sky130_fd_sc_hd__or2b_2 c559(
.A(net338),
.B_N(net852),
.X(net449)
);

sky130_fd_sc_hd__clkinv_4 c560(
.A(out15),
.Y(net450)
);

sky130_fd_sc_hd__and3b_4 c561(
.A_N(net319),
.B(net333),
.C(net837),
.X(net451)
);

sky130_fd_sc_hd__nand2b_1 c562(
.A_N(net437),
.B(net442),
.Y(net452)
);

sky130_fd_sc_hd__inv_12 c563(
.A(net801),
.Y(net453)
);

sky130_fd_sc_hd__buf_12 c564(
.A(net807),
.X(net454)
);

sky130_fd_sc_hd__and3_4 c565(
.A(net452),
.B(net449),
.C(net433),
.X(net455)
);

sky130_fd_sc_hd__o211a_1 c566(
.A1(net448),
.A2(net455),
.B1(net433),
.C1(net861),
.X(net456)
);

sky130_fd_sc_hd__clkbuf_16 c567(
.A(net801),
.X(net457)
);

sky130_fd_sc_hd__or3_1 c568(
.A(net433),
.B(net453),
.C(net457),
.X(net458)
);

sky130_fd_sc_hd__sdfbbn_1 c569(
.D(net316),
.RESET_B(net447),
.SCD(net458),
.SCE(net445),
.SET_B(net457),
.CLK_N(clk),
.Q(net460),
.Q_N(net459)
);

sky130_fd_sc_hd__o211ai_2 c570(
.A1(net457),
.A2(net455),
.B1(net459),
.C1(net752),
.Y(net461)
);

sky130_fd_sc_hd__sdfbbn_2 c571(
.D(net455),
.RESET_B(net454),
.SCD(net427),
.SCE(net457),
.SET_B(net752),
.CLK_N(clk),
.Q(net463),
.Q_N(net462)
);

sky130_fd_sc_hd__nand3_4 c572(
.A(net460),
.B(net429),
.C(net333),
.Y(net464)
);

sky130_fd_sc_hd__o221ai_4 c573(
.A1(in47),
.A2(net460),
.B1(net429),
.B2(net417),
.C1(net362),
.Y(net465)
);

sky130_fd_sc_hd__o221a_2 c574(
.A1(net362),
.A2(net429),
.B1(out19),
.B2(net94),
.C1(net333),
.X(net466)
);

sky130_fd_sc_hd__clkinv_1 c575(
.A(net786),
.Y(net467)
);

sky130_fd_sc_hd__buf_1 c576(
.A(net786),
.X(net468)
);

sky130_fd_sc_hd__o221a_2 c577(
.A1(net460),
.A2(net468),
.B1(net711),
.B2(net799),
.C1(net857),
.X(net469)
);

sky130_fd_sc_hd__o221a_2 c578(
.A1(net308),
.A2(net318),
.B1(net446),
.B2(net857),
.C1(net862),
.X(net470)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c579(
.A(net800),
.X(net471)
);

sky130_fd_sc_hd__mux4_2 c580(
.A0(net469),
.A1(net72),
.A2(net445),
.A3(net417),
.S0(out19),
.S1(net333),
.X(net472)
);

sky130_fd_sc_hd__clkinv_8 c581(
.A(net776),
.Y(net473)
);

sky130_fd_sc_hd__mux4_2 c582(
.A0(net473),
.A1(net417),
.A2(net469),
.A3(in3),
.S0(in47),
.S1(net862),
.X(net474)
);

sky130_fd_sc_hd__mux4_4 c583(
.A0(net470),
.A1(net94),
.A2(net429),
.A3(net728),
.S0(net863),
.S1(net865),
.X(net475)
);

sky130_fd_sc_hd__o221ai_1 c584(
.A1(in56),
.A2(net318),
.B1(net446),
.B2(net857),
.C1(net865),
.Y(net476)
);

sky130_fd_sc_hd__mux4_1 c585(
.A0(net469),
.A1(net333),
.A2(net476),
.A3(net857),
.S0(net862),
.S1(net865),
.X(net477)
);

sky130_fd_sc_hd__mux4_1 c586(
.A0(net94),
.A1(in35),
.A2(net463),
.A3(net800),
.S0(net864),
.S1(net865),
.X(net478)
);

sky130_fd_sc_hd__sdfbbp_1 c587(
.D(net467),
.RESET_B(net362),
.SCD(net476),
.SCE(net857),
.SET_B(net865),
.CLK(clk),
.Q(net480),
.Q_N(net479)
);

sky130_fd_sc_hd__mux4_1 c588(
.A0(net478),
.A1(net480),
.A2(net125),
.A3(net254),
.S0(net459),
.S1(net457),
.X(net481)
);

sky130_fd_sc_hd__mux4_4 c589(
.A0(net468),
.A1(net478),
.A2(net94),
.A3(net481),
.S0(out3),
.S1(net865),
.X(net482)
);

sky130_fd_sc_hd__mux4_1 c590(
.A0(net429),
.A1(net481),
.A2(net468),
.A3(net476),
.S0(net799),
.S1(net867),
.X(net483)
);

sky130_fd_sc_hd__mux4_4 c591(
.A0(net446),
.A1(net480),
.A2(out2),
.A3(net468),
.S0(net457),
.S1(net862),
.X(net484)
);

sky130_fd_sc_hd__mux4_4 c592(
.A0(net247),
.A1(net478),
.A2(net479),
.A3(net429),
.S0(net800),
.S1(net866),
.X(net485)
);

sky130_fd_sc_hd__mux4_2 c593(
.A0(net471),
.A1(net463),
.A2(net485),
.A3(net417),
.S0(net468),
.S1(net712),
.X(net486)
);

sky130_fd_sc_hd__clkbuf_2 c594(
.A(net814),
.X(net487)
);

sky130_fd_sc_hd__o211a_2 c595(
.A1(net422),
.A2(net94),
.B1(net457),
.C1(net841),
.X(net488)
);

sky130_fd_sc_hd__o221a_2 c596(
.A1(net386),
.A2(net260),
.B1(net5),
.B2(net207),
.C1(net484),
.X(net489)
);

sky130_fd_sc_hd__mux4_4 c597(
.A0(net264),
.A1(out19),
.A2(net353),
.A3(in32),
.S0(net464),
.S1(net94),
.X(net490)
);

sky130_fd_sc_hd__o221a_2 c598(
.A1(in32),
.A2(net376),
.B1(net476),
.B2(net94),
.C1(net832),
.X(net491)
);

sky130_fd_sc_hd__o221ai_1 c599(
.A1(net207),
.A2(net8),
.B1(net319),
.B2(net840),
.C1(net869),
.Y(net492)
);

sky130_fd_sc_hd__mux4_4 c600(
.A0(net422),
.A1(net283),
.A2(net372),
.A3(net712),
.S0(out4),
.S1(net868),
.X(net493)
);

sky130_fd_sc_hd__sdfbbn_1 c601(
.D(net484),
.RESET_B(net457),
.SCD(net476),
.SCE(net94),
.SET_B(net5),
.CLK_N(clk),
.Q(net495),
.Q_N(net494)
);

sky130_fd_sc_hd__o221a_4 c602(
.A1(net492),
.A2(net142),
.B1(net457),
.B2(out38),
.C1(net868),
.X(net496)
);

sky130_fd_sc_hd__sdfbbn_2 c603(
.D(net5),
.RESET_B(out19),
.SCD(net422),
.SCE(net72),
.SET_B(net869),
.CLK_N(clk),
.Q(net498),
.Q_N(net497)
);

sky130_fd_sc_hd__o221a_2 c604(
.A1(net476),
.A2(net277),
.B1(net281),
.B2(net496),
.C1(out17),
.X(net499)
);

sky130_fd_sc_hd__o221ai_4 c605(
.A1(net487),
.A2(net8),
.B1(out3),
.B2(net866),
.C1(out17),
.Y(net500)
);

sky130_fd_sc_hd__o221a_2 c606(
.A1(net487),
.A2(net498),
.B1(net494),
.B2(out19),
.C1(out8),
.X(net501)
);

sky130_fd_sc_hd__o221a_1 c607(
.A1(net246),
.A2(net500),
.B1(net386),
.B2(net320),
.C1(net832),
.X(net502)
);

sky130_fd_sc_hd__or3b_1 c608(
.A(net497),
.B(out15),
.C_N(out9),
.X(net503)
);

sky130_fd_sc_hd__o221ai_1 c609(
.A1(net385),
.A2(net387),
.B1(net487),
.B2(net503),
.C1(net869),
.Y(net504)
);

sky130_fd_sc_hd__mux4_4 c610(
.A0(net488),
.A1(net503),
.A2(net497),
.A3(net504),
.S0(net457),
.S1(net811),
.X(net505)
);

sky130_fd_sc_hd__mux4_2 c611(
.A0(net495),
.A1(net503),
.A2(net284),
.A3(net504),
.S0(net72),
.S1(net92),
.X(net506)
);

sky130_fd_sc_hd__mux4_4 c612(
.A0(net387),
.A1(net495),
.A2(net504),
.A3(net503),
.S0(net811),
.S1(net870),
.X(net507)
);

sky130_fd_sc_hd__clkbuf_1 c613(
.A(net814),
.X(net508)
);

sky130_fd_sc_hd__mux4_2 c614(
.A0(net496),
.A1(net503),
.A2(net142),
.A3(net353),
.S0(net494),
.S1(net870),
.X(net509)
);

sky130_fd_sc_hd__mux4_2 c615(
.A0(net509),
.A1(net495),
.A2(net488),
.A3(net503),
.S0(net508),
.S1(out11),
.X(net510)
);

sky130_fd_sc_hd__mux4_1 c616(
.A0(net262),
.A1(net34),
.A2(out19),
.A3(net846),
.S0(out3),
.S1(net873),
.X(net511)
);

sky130_fd_sc_hd__mux4_4 c617(
.A0(net169),
.A1(out2),
.A2(net320),
.A3(net858),
.S0(net860),
.S1(net868),
.X(net512)
);

sky130_fd_sc_hd__mux4_1 c618(
.A0(net281),
.A1(net94),
.A2(net72),
.A3(in32),
.S0(net844),
.S1(net867),
.X(net513)
);

sky130_fd_sc_hd__mux4_4 c619(
.A0(net498),
.A1(out7),
.A2(net162),
.A3(net464),
.S0(net835),
.S1(net860),
.X(net514)
);

sky130_fd_sc_hd__mux4_2 c620(
.A0(net303),
.A1(net513),
.A2(net498),
.A3(net457),
.S0(net860),
.S1(net875),
.X(net515)
);

sky130_fd_sc_hd__mux4_4 c621(
.A0(net162),
.A1(in31),
.A2(out10),
.A3(net257),
.S0(net840),
.S1(out3),
.X(net516)
);

sky130_fd_sc_hd__mux4_1 c622(
.A0(net34),
.A1(net303),
.A2(net780),
.A3(out0),
.S0(net843),
.S1(net860),
.X(net517)
);

sky130_fd_sc_hd__mux4_2 c623(
.A0(net320),
.A1(net513),
.A2(net464),
.A3(out11),
.S0(out4),
.S1(net868),
.X(net518)
);

sky130_fd_sc_hd__mux4_4 c624(
.A0(in16),
.A1(net372),
.A2(out7),
.A3(net94),
.S0(net422),
.S1(net870),
.X(net519)
);

sky130_fd_sc_hd__mux4_4 c625(
.A0(net94),
.A1(net516),
.A2(out16),
.A3(net389),
.S0(net840),
.S1(net858),
.X(net520)
);

sky130_fd_sc_hd__mux4_2 c626(
.A0(net513),
.A1(net389),
.A2(net796),
.A3(net825),
.S0(net858),
.S1(net874),
.X(net521)
);

sky130_fd_sc_hd__mux4_2 c627(
.A0(in35),
.A1(net487),
.A2(net257),
.A3(net72),
.S0(out2),
.S1(out25),
.X(net522)
);

sky130_fd_sc_hd__mux4_1 c628(
.A0(net522),
.A1(net42),
.A2(out1),
.A3(net457),
.S0(net844),
.S1(out38),
.X(net523)
);

sky130_fd_sc_hd__mux4_1 c629(
.A0(net521),
.A1(net257),
.A2(net513),
.A3(net162),
.S0(net816),
.S1(net860),
.X(net524)
);

sky130_fd_sc_hd__mux4_1 c630(
.A0(net34),
.A1(net521),
.A2(net169),
.A3(net825),
.S0(net860),
.S1(out20),
.X(net525)
);

sky130_fd_sc_hd__mux4_2 c631(
.A0(net422),
.A1(net293),
.A2(net513),
.A3(out16),
.S0(net780),
.S1(net858),
.X(out13)
);

sky130_fd_sc_hd__mux4_2 c632(
.A0(out13),
.A1(net464),
.A2(net513),
.A3(net508),
.S0(net803),
.S1(net815),
.X(net526)
);

sky130_fd_sc_hd__mux4_1 c633(
.A0(net457),
.A1(net521),
.A2(net422),
.A3(net513),
.S0(net845),
.S1(net867),
.X(net527)
);

sky130_fd_sc_hd__mux4_1 c634(
.A0(net257),
.A1(net42),
.A2(net835),
.A3(net860),
.S0(net867),
.S1(net876),
.X(net528)
);

sky130_fd_sc_hd__mux4_1 c635(
.A0(net528),
.A1(net457),
.A2(net169),
.A3(net422),
.S0(out17),
.S1(net876),
.X(net529)
);

sky130_fd_sc_hd__mux4_1 c636(
.A0(out10),
.A1(net528),
.A2(net41),
.A3(net816),
.S0(out38),
.S1(net877),
.X(net530)
);

sky130_fd_sc_hd__mux4_4 c637(
.A0(net530),
.A1(net284),
.A2(in29),
.A3(out19),
.S0(net840),
.S1(net877),
.X(net531)
);

sky130_fd_sc_hd__or2b_1 c660(
.A(net81),
.B_N(net434),
.X(net532)
);

sky130_fd_sc_hd__buf_6 c661(
.A(net806),
.X(net533)
);

sky130_fd_sc_hd__clkinv_8 c662(
.A(net646),
.Y(net534)
);

sky130_fd_sc_hd__buf_16 c663(
.A(net645),
.X(net535)
);

sky130_fd_sc_hd__nand3_1 c664(
.A(net432),
.B(net215),
.C(net81),
.Y(net536)
);

sky130_fd_sc_hd__inv_6 c665(
.A(net817),
.Y(net537)
);

sky130_fd_sc_hd__sdfrtp_1 c666(
.D(net424),
.RESET_B(net532),
.SCD(net78),
.SCE(net535),
.CLK(clk),
.Q(net538)
);

sky130_fd_sc_hd__inv_12 c667(
.A(net817),
.Y(net539)
);

sky130_fd_sc_hd__clkinv_2 c668(
.A(net761),
.Y(net540)
);

sky130_fd_sc_hd__nand2b_1 c669(
.A_N(net86),
.B(net848),
.Y(net541)
);

sky130_fd_sc_hd__or2_1 c670(
.A(net540),
.B(net204),
.X(net542)
);

sky130_fd_sc_hd__or2_1 c671(
.A(net416),
.B(net542),
.X(net543)
);

sky130_fd_sc_hd__mux4_1 c672(
.A0(net536),
.A1(net541),
.A2(net317),
.A3(net534),
.S0(net539),
.S1(net309),
.X(net544)
);

sky130_fd_sc_hd__buf_6 c673(
.A(net792),
.X(net545)
);

sky130_fd_sc_hd__nand2b_1 c674(
.A_N(net541),
.B(net545),
.Y(net546)
);

sky130_fd_sc_hd__nand2_1 c675(
.A(net317),
.B(net204),
.Y(net547)
);

sky130_fd_sc_hd__mux4_4 c676(
.A0(net533),
.A1(net543),
.A2(net539),
.A3(net540),
.S0(net545),
.S1(net879),
.X(net548)
);

sky130_fd_sc_hd__clkinv_8 c677(
.A(net761),
.Y(net549)
);

sky130_fd_sc_hd__mux4_2 c678(
.A0(net208),
.A1(net542),
.A2(net549),
.A3(net548),
.S0(net545),
.S1(net538),
.X(net550)
);

sky130_fd_sc_hd__or3_2 c679(
.A(net545),
.B(net543),
.C(net772),
.X(net551)
);

sky130_fd_sc_hd__mux4_1 c680(
.A0(net549),
.A1(net551),
.A2(net317),
.A3(net548),
.S0(net532),
.S1(net543),
.X(net552)
);

sky130_fd_sc_hd__sdfbbp_1 c681(
.D(net438),
.RESET_B(net548),
.SCD(net551),
.SCE(net324),
.SET_B(net772),
.CLK(clk),
.Q(net554),
.Q_N(net553)
);

sky130_fd_sc_hd__nand3b_2 c682(
.A_N(net537),
.B(net547),
.C(net72),
.Y(net555)
);

sky130_fd_sc_hd__sdfrtp_2 c683(
.D(net548),
.RESET_B(net538),
.SCD(net457),
.SCE(net879),
.CLK(clk),
.Q(net556)
);

sky130_fd_sc_hd__o211a_4 c684(
.A1(net554),
.A2(net535),
.B1(in32),
.C1(net879),
.X(net557)
);

sky130_fd_sc_hd__nand3_4 c685(
.A(net557),
.B(net537),
.C(net556),
.Y(net558)
);

sky130_fd_sc_hd__o211a_1 c686(
.A1(net558),
.A2(net547),
.B1(net548),
.C1(net457),
.X(net559)
);

sky130_fd_sc_hd__sdfbbn_1 c687(
.D(net543),
.RESET_B(net558),
.SCD(net78),
.SCE(net555),
.SET_B(net553),
.CLK_N(clk),
.Q(net561),
.Q_N(net560)
);

sky130_fd_sc_hd__sdfrtp_4 c688(
.D(net555),
.RESET_B(net545),
.SCD(net557),
.SCE(net457),
.CLK(clk),
.Q(net562)
);

sky130_fd_sc_hd__mux4_2 c689(
.A0(net547),
.A1(net555),
.A2(net556),
.A3(net543),
.S0(net561),
.S1(net535),
.X(net563)
);

sky130_fd_sc_hd__sdfbbn_2 c690(
.D(net200),
.RESET_B(net558),
.SCD(in32),
.SCE(net557),
.SET_B(net556),
.CLK_N(clk),
.Q(net565),
.Q_N(net564)
);

sky130_fd_sc_hd__mux4_4 c691(
.A0(net85),
.A1(net558),
.A2(net545),
.A3(net557),
.S0(net458),
.S1(net880),
.X(net566)
);

sky130_fd_sc_hd__o221a_4 c692(
.A1(net454),
.A2(net554),
.B1(net564),
.B2(net458),
.C1(net457),
.X(net567)
);

sky130_fd_sc_hd__o221ai_1 c693(
.A1(net567),
.A2(net448),
.B1(net562),
.B2(net537),
.C1(net457),
.Y(net568)
);

sky130_fd_sc_hd__mux4_4 c694(
.A0(net561),
.A1(net538),
.A2(in16),
.A3(net556),
.S0(net85),
.S1(net457),
.X(net569)
);

sky130_fd_sc_hd__inv_12 c695(
.A(out15),
.Y(net570)
);

sky130_fd_sc_hd__mux4_2 c696(
.A0(net569),
.A1(in31),
.A2(net553),
.A3(net564),
.S0(net454),
.S1(net560),
.X(net571)
);

sky130_fd_sc_hd__and3b_1 c697(
.A_N(net538),
.B(net556),
.C(net458),
.X(net572)
);

sky130_fd_sc_hd__o221a_2 c698(
.A1(net570),
.A2(net548),
.B1(net572),
.B2(net560),
.C1(net535),
.X(net573)
);

sky130_fd_sc_hd__mux4_2 c699(
.A0(net566),
.A1(net458),
.A2(net556),
.A3(net535),
.S0(net564),
.S1(net883),
.X(net574)
);

sky130_fd_sc_hd__mux4_2 c700(
.A0(net572),
.A1(net557),
.A2(net556),
.A3(net454),
.S0(net457),
.S1(net795),
.X(net575)
);

sky130_fd_sc_hd__sdfbbp_1 c701(
.D(net556),
.RESET_B(net545),
.SCD(net532),
.SCE(net572),
.SET_B(net457),
.CLK(clk),
.Q(net577),
.Q_N(net576)
);

sky130_fd_sc_hd__mux4_2 c702(
.A0(net575),
.A1(net577),
.A2(net558),
.A3(net538),
.S0(net572),
.S1(net761),
.X(net578)
);

sky130_fd_sc_hd__mux4_1 c703(
.A0(net78),
.A1(net562),
.A2(net572),
.A3(net577),
.S0(net564),
.S1(net883),
.X(net579)
);

sky130_fd_sc_hd__sdfbbn_1 c704(
.D(net485),
.RESET_B(net125),
.SCD(net577),
.SCE(net562),
.SET_B(net882),
.CLK_N(clk),
.Q(net581),
.Q_N(net580)
);

sky130_fd_sc_hd__o221a_4 c705(
.A1(net318),
.A2(net125),
.B1(net565),
.B2(net485),
.C1(net535),
.X(net582)
);

sky130_fd_sc_hd__mux4_4 c706(
.A0(net485),
.A1(net535),
.A2(net581),
.A3(net458),
.S0(out43),
.S1(net864),
.X(net583)
);

sky130_fd_sc_hd__sdfbbn_2 c707(
.D(net577),
.RESET_B(net546),
.SCD(net458),
.SCE(net580),
.SET_B(net880),
.CLK_N(clk),
.Q(net585),
.Q_N(net584)
);

sky130_fd_sc_hd__o211a_2 c708(
.A1(net535),
.A2(net125),
.B1(in3),
.C1(net864),
.X(net586)
);

sky130_fd_sc_hd__o221ai_4 c709(
.A1(net565),
.A2(in29),
.B1(net580),
.B2(net94),
.C1(net883),
.Y(net587)
);

sky130_fd_sc_hd__o221ai_1 c710(
.A1(net585),
.A2(in3),
.B1(in16),
.B2(net94),
.C1(net817),
.Y(net588)
);

sky130_fd_sc_hd__o221a_4 c711(
.A1(net215),
.A2(net535),
.B1(net576),
.B2(net866),
.C1(net882),
.X(net589)
);

sky130_fd_sc_hd__mux4_1 c712(
.A0(net546),
.A1(net589),
.A2(net577),
.A3(net584),
.S0(net457),
.S1(net728),
.X(net590)
);

sky130_fd_sc_hd__o211ai_4 c713(
.A1(net585),
.A2(net125),
.B1(net589),
.C1(net883),
.Y(net591)
);

sky130_fd_sc_hd__mux4_1 c714(
.A0(net589),
.A1(net579),
.A2(net72),
.A3(net580),
.S0(net532),
.S1(net882),
.X(net592)
);

sky130_fd_sc_hd__o221ai_4 c715(
.A1(net576),
.A2(net761),
.B1(net817),
.B2(net866),
.C1(net884),
.Y(net593)
);

sky130_fd_sc_hd__sdfbbp_1 c716(
.D(net593),
.RESET_B(net485),
.SCD(net535),
.SCE(net580),
.SET_B(net863),
.CLK(clk),
.Q(net595),
.Q_N(net594)
);

sky130_fd_sc_hd__o221a_2 c717(
.A1(net458),
.A2(net584),
.B1(net565),
.B2(net588),
.C1(net576),
.X(net596)
);

sky130_fd_sc_hd__sdfbbn_1 c718(
.D(net532),
.RESET_B(net595),
.SCD(net565),
.SCE(net863),
.SET_B(net881),
.CLK_N(clk),
.Q(net598),
.Q_N(net597)
);

sky130_fd_sc_hd__mux4_1 c719(
.A0(net586),
.A1(net125),
.A2(net576),
.A3(net458),
.S0(net588),
.S1(net885),
.X(net599)
);

sky130_fd_sc_hd__mux4_4 c720(
.A0(net596),
.A1(net599),
.A2(net458),
.A3(net795),
.S0(net882),
.S1(net885),
.X(net600)
);

sky130_fd_sc_hd__o221ai_1 c721(
.A1(net586),
.A2(net594),
.B1(net867),
.B2(net883),
.C1(net886),
.Y(net601)
);

sky130_fd_sc_hd__o221a_1 c722(
.A1(net581),
.A2(net485),
.B1(net601),
.B2(net125),
.C1(net758),
.X(net602)
);

sky130_fd_sc_hd__mux4_4 c723(
.A0(net599),
.A1(net581),
.A2(in16),
.A3(net758),
.S0(net885),
.S1(net886),
.X(net603)
);

sky130_fd_sc_hd__mux4_2 c724(
.A0(net601),
.A1(net599),
.A2(net589),
.A3(net597),
.S0(in31),
.S1(net795),
.X(net604)
);

sky130_fd_sc_hd__mux4_1 c725(
.A0(net587),
.A1(net596),
.A2(net565),
.A3(net758),
.S0(net795),
.S1(net886),
.X(net605)
);

sky130_fd_sc_hd__mux4_4 c726(
.A0(net581),
.A1(net309),
.A2(in31),
.A3(net866),
.S0(net871),
.S1(net873),
.X(net606)
);

sky130_fd_sc_hd__o221ai_4 c727(
.A1(net142),
.A2(net588),
.B1(net562),
.B2(net551),
.C1(net886),
.Y(net607)
);

sky130_fd_sc_hd__mux4_2 c728(
.A0(net254),
.A1(net376),
.A2(net551),
.A3(net8),
.S0(net791),
.S1(net884),
.X(net608)
);

sky130_fd_sc_hd__mux4_4 c729(
.A0(net309),
.A1(net551),
.A2(net580),
.A3(net8),
.S0(net866),
.S1(net871),
.X(net609)
);

sky130_fd_sc_hd__mux4_4 c730(
.A0(net551),
.A1(net598),
.A2(net562),
.A3(net799),
.S0(net832),
.S1(out4),
.X(net610)
);

sky130_fd_sc_hd__mux4_4 c731(
.A0(net599),
.A1(net284),
.A2(net562),
.A3(in3),
.S0(net868),
.S1(net888),
.X(net611)
);

sky130_fd_sc_hd__mux4_2 c732(
.A0(net382),
.A1(in16),
.A2(net283),
.A3(net791),
.S0(net798),
.S1(net887),
.X(net612)
);

sky130_fd_sc_hd__mux4_2 c733(
.A0(net374),
.A1(net595),
.A2(net8),
.A3(net309),
.S0(net457),
.S1(net866),
.X(net613)
);

sky130_fd_sc_hd__mux4_2 c734(
.A0(net612),
.A1(net374),
.A2(net283),
.A3(in3),
.S0(net885),
.S1(net888),
.X(net614)
);

sky130_fd_sc_hd__mux4_1 c735(
.A0(net601),
.A1(net546),
.A2(net581),
.A3(in32),
.S0(out4),
.S1(net881),
.X(net615)
);

sky130_fd_sc_hd__o221a_2 c736(
.A1(net581),
.A2(net383),
.B1(net612),
.B2(net798),
.C1(net811),
.X(net616)
);

sky130_fd_sc_hd__mux4_4 c737(
.A0(net616),
.A1(net376),
.A2(net254),
.A3(net770),
.S0(net821),
.S1(net881),
.X(net617)
);

sky130_fd_sc_hd__o221ai_2 c738(
.A1(net8),
.A2(in3),
.B1(net562),
.B2(net551),
.C1(net811),
.Y(net618)
);

sky130_fd_sc_hd__mux4_2 c739(
.A0(net387),
.A1(net464),
.A2(net617),
.A3(net142),
.S0(net803),
.S1(net884),
.X(net619)
);

sky130_fd_sc_hd__mux4_1 c740(
.A0(net383),
.A1(net125),
.A2(net309),
.A3(net616),
.S0(net94),
.S1(net868),
.X(net620)
);

sky130_fd_sc_hd__mux4_4 c741(
.A0(net617),
.A1(net824),
.A2(out11),
.A3(net832),
.S0(net868),
.S1(net890),
.X(net621)
);

sky130_fd_sc_hd__o221ai_4 c742(
.A1(net562),
.A2(net601),
.B1(net374),
.B2(net888),
.C1(net891),
.Y(net622)
);

sky130_fd_sc_hd__o221ai_4 c743(
.A1(net617),
.A2(net309),
.B1(net822),
.B2(net880),
.C1(net890),
.Y(net623)
);

sky130_fd_sc_hd__o221a_2 c744(
.A1(net617),
.A2(net309),
.B1(net616),
.B2(net822),
.C1(net881),
.X(net624)
);

sky130_fd_sc_hd__mux4_4 c745(
.A0(net142),
.A1(net612),
.A2(net617),
.A3(net546),
.S0(net821),
.S1(net889),
.X(net625)
);

sky130_fd_sc_hd__mux4_1 c746(
.A0(net616),
.A1(in29),
.A2(net464),
.A3(net770),
.S0(net796),
.S1(net890),
.X(net626)
);

sky130_fd_sc_hd__mux4_4 c747(
.A0(net617),
.A1(net508),
.A2(net387),
.A3(net785),
.S0(net880),
.S1(net892),
.X(net627)
);

sky130_fd_sc_hd__mux4_4 c748(
.A0(net72),
.A1(in32),
.A2(net866),
.A3(net873),
.S0(net875),
.S1(net894),
.X(net628)
);

sky130_fd_sc_hd__mux4_1 c749(
.A0(net284),
.A1(in31),
.A2(out4),
.A3(net874),
.S0(net889),
.S1(net891),
.X(net629)
);

sky130_fd_sc_hd__mux4_4 c750(
.A0(net546),
.A1(net867),
.A2(net871),
.A3(net872),
.S0(net891),
.S1(net893),
.X(net630)
);

sky130_fd_sc_hd__mux4_4 c751(
.A0(in32),
.A1(net799),
.A2(net874),
.A3(net878),
.S0(net892),
.S1(net895),
.X(net631)
);

sky130_fd_sc_hd__mux4_2 c752(
.A0(net588),
.A1(out4),
.A2(net878),
.A3(net889),
.S0(net891),
.S1(net895),
.X(net632)
);

sky130_fd_sc_hd__mux4_2 c753(
.A0(net628),
.A1(net632),
.A2(net588),
.A3(net867),
.S0(net874),
.S1(net893),
.X(net633)
);

sky130_fd_sc_hd__mux4_4 c754(
.A0(net631),
.A1(in31),
.A2(net781),
.A3(out4),
.S0(net875),
.S1(net894),
.X(net634)
);

sky130_fd_sc_hd__mux4_2 c755(
.A0(net588),
.A1(net516),
.A2(net508),
.A3(net796),
.S0(net868),
.S1(net894),
.X(net635)
);

sky130_fd_sc_hd__mux4_4 c756(
.A0(net72),
.A1(net283),
.A2(net796),
.A3(net866),
.S0(net878),
.S1(net896),
.X(net636)
);

sky130_fd_sc_hd__mux4_4 c757(
.A0(net464),
.A1(in16),
.A2(net546),
.A3(net781),
.S0(net887),
.S1(net896),
.X(net637)
);

sky130_fd_sc_hd__mux4_2 c758(
.A0(net629),
.A1(net866),
.A2(net868),
.A3(net894),
.S0(net896),
.S1(net897),
.X(net638)
);

sky130_fd_sc_hd__mux4_2 c759(
.A0(net508),
.A1(net464),
.A2(net887),
.A3(net889),
.S0(net895),
.S1(net896),
.X(net639)
);

sky130_fd_sc_hd__mux4_1 c760(
.A0(net636),
.A1(net546),
.A2(net872),
.A3(net887),
.S0(net896),
.S1(net897),
.X(net640)
);

sky130_fd_sc_hd__mux4_2 c761(
.A0(net598),
.A1(net824),
.A2(net871),
.A3(net889),
.S0(net896),
.S1(net897),
.X(net641)
);

sky130_fd_sc_hd__mux4_4 c762(
.A0(net634),
.A1(net284),
.A2(net546),
.A3(net867),
.S0(net893),
.S1(net896),
.X(net642)
);

sky130_fd_sc_hd__mux4_1 c763(
.A0(net641),
.A1(net508),
.A2(net803),
.A3(net875),
.S0(net884),
.S1(net896),
.X(net643)
);

sky130_fd_sc_hd__mux4_2 c764(
.A0(net638),
.A1(net643),
.A2(net508),
.A3(net803),
.S0(net875),
.S1(net895)
);

sky130_fd_sc_hd__mux4_1 merge765(
.A0(net332),
.A1(net200),
.A2(net308),
.A3(net330),
.S0(net336),
.S1(net333),
.X(net644)
);

sky130_fd_sc_hd__sdfsbp_1 merge766(
.D(net430),
.SCD(net438),
.SCE(net204),
.SET_B(net532),
.CLK(clk),
.Q(net646),
.Q_N(net645)
);

sky130_fd_sc_hd__o221ai_2 merge767(
.A1(in38),
.A2(net80),
.B1(net102),
.B2(net95),
.C1(net94),
.Y(net647)
);

sky130_fd_sc_hd__o211ai_1 merge768(
.A1(net103),
.A2(net122),
.B1(net124),
.C1(net121),
.Y(net648)
);

sky130_fd_sc_hd__o211a_4 merge769(
.A1(net76),
.A2(net72),
.B1(in19),
.C1(net80),
.X(net649)
);

sky130_fd_sc_hd__o211a_1 merge770(
.A1(net200),
.A2(net81),
.B1(net205),
.C1(net203),
.X(net650)
);

sky130_fd_sc_hd__o211ai_1 merge771(
.A1(net0),
.A2(out56),
.B1(net234),
.C1(net267),
.Y(net651)
);

sky130_fd_sc_hd__o211ai_1 merge772(
.A1(net223),
.A2(net224),
.B1(net205),
.C1(net233),
.Y(net652)
);

sky130_fd_sc_hd__o221a_1 merge773(
.A1(net333),
.A2(net445),
.B1(net417),
.B2(net362),
.C1(net861),
.X(net653)
);

sky130_fd_sc_hd__inv_6 merge774(
.A(net777),
.Y(net654)
);

sky130_fd_sc_hd__o221ai_2 merge775(
.A1(net239),
.A2(net234),
.B1(net128),
.B2(net237),
.C1(net130),
.Y(net655)
);

sky130_fd_sc_hd__mux4_2 merge776(
.A0(net319),
.A1(net476),
.A2(net246),
.A3(net504),
.S0(net494),
.S1(net503),
.X(net656)
);

sky130_fd_sc_hd__o211a_1 merge777(
.A1(in36),
.A2(out30),
.B1(net26),
.C1(net25),
.X(net657)
);

sky130_fd_sc_hd__o211ai_1 merge778(
.A1(net347),
.A2(net427),
.B1(net849),
.C1(net851),
.Y(net658)
);

sky130_fd_sc_hd__o211ai_2 merge779(
.A1(net91),
.A2(net315),
.B1(net417),
.C1(net316),
.Y(net659)
);

sky130_fd_sc_hd__o211ai_1 merge780(
.A1(net90),
.A2(in0),
.B1(net308),
.C1(net309),
.Y(net660)
);

sky130_fd_sc_hd__clkinv_4 merge781(
.A(net793),
.Y(net661)
);

sky130_fd_sc_hd__mux4_2 merge782(
.A0(net18),
.A1(out56),
.A2(net55),
.A3(in21),
.S0(net160),
.S1(net779),
.X(net662)
);

sky130_fd_sc_hd__mux4_1 merge783(
.A0(net356),
.A1(net363),
.A2(net277),
.A3(net350),
.S0(net281),
.S1(net835),
.X(net663)
);

sky130_fd_sc_hd__o211a_1 merge784(
.A1(net152),
.A2(out52),
.B1(net167),
.C1(net729),
.X(net664)
);

sky130_fd_sc_hd__mux4_1 merge785(
.A0(net354),
.A1(out33),
.A2(net351),
.A3(net357),
.S0(net333),
.S1(net839),
.X(net665)
);

sky130_fd_sc_hd__mux4_1 merge786(
.A0(net278),
.A1(net34),
.A2(net45),
.A3(net178),
.S0(out10),
.S1(out58),
.X(net666)
);

sky130_fd_sc_hd__o211a_2 merge787(
.A1(net111),
.A2(net146),
.B1(out55),
.C1(net820),
.X(net667)
);

sky130_fd_sc_hd__o221ai_2 merge788(
.A1(net16),
.A2(net0),
.B1(net224),
.B2(net21),
.C1(out52),
.Y(net668)
);

sky130_fd_sc_hd__clkinv_4 merge789(
.A(net810),
.Y(net669)
);

sky130_fd_sc_hd__mux4_4 merge790(
.A0(net568),
.A1(net562),
.A2(net454),
.A3(net442),
.S0(net445),
.S1(out19),
.X(net670)
);

sky130_fd_sc_hd__o211ai_4 merge791(
.A1(net315),
.A2(net427),
.B1(net76),
.C1(net309),
.Y(net671)
);

sky130_fd_sc_hd__mux4_2 merge792(
.A0(net372),
.A1(net5),
.A2(out36),
.A3(net175),
.S0(net150),
.S1(net41),
.X(net672)
);

sky130_fd_sc_hd__o211ai_4 merge793(
.A1(net434),
.A2(net309),
.B1(net438),
.C1(net424),
.Y(net673)
);

sky130_fd_sc_hd__mux4_4 merge794(
.A0(net297),
.A1(net273),
.A2(net34),
.A3(net127),
.S0(out52),
.S1(net729),
.X(net674)
);

sky130_fd_sc_hd__mux4_4 merge795(
.A0(in54),
.A1(out55),
.A2(out6),
.A3(net294),
.S0(net290),
.S1(out1),
.X(net675)
);

sky130_fd_sc_hd__o211a_1 merge796(
.A1(net213),
.A2(net209),
.B1(net238),
.C1(net234),
.X(net676)
);

sky130_fd_sc_hd__o211a_2 merge797(
.A1(net315),
.A2(net309),
.B1(net320),
.C1(net312),
.X(net677)
);

sky130_fd_sc_hd__o211ai_4 merge798(
.A1(net206),
.A2(net203),
.B1(net80),
.C1(in8),
.Y(net678)
);

sky130_fd_sc_hd__o211ai_2 merge799(
.A1(net237),
.A2(net73),
.B1(net200),
.C1(net812),
.Y(net679)
);

sky130_fd_sc_hd__o221ai_1 merge800(
.A1(net539),
.A2(net536),
.B1(net534),
.B2(net548),
.C1(net547),
.Y(net680)
);

sky130_fd_sc_hd__mux4_2 merge801(
.A0(net13),
.A1(net16),
.A2(net8),
.A3(net95),
.S0(net103),
.S1(net102),
.X(net681)
);

sky130_fd_sc_hd__mux4_2 merge802(
.A0(net245),
.A1(net464),
.A2(net429),
.A3(net361),
.S0(net71),
.S1(out38),
.X(net682)
);

sky130_fd_sc_hd__mux4_4 merge803(
.A0(net119),
.A1(net361),
.A2(net353),
.A3(net88),
.S0(net124),
.S1(net114),
.X(net683)
);

sky130_fd_sc_hd__mux4_2 merge804(
.A0(net110),
.A1(net106),
.A2(net96),
.A3(net273),
.S0(net213),
.S1(net818),
.X(net684)
);

sky130_fd_sc_hd__o211ai_4 merge805(
.A1(net38),
.A2(out30),
.B1(net65),
.C1(net826),
.Y(net685)
);

sky130_fd_sc_hd__mux4_1 merge806(
.A0(net30),
.A1(net26),
.A2(net11),
.A3(net182),
.S0(net180),
.S1(out57),
.X(net686)
);

sky130_fd_sc_hd__mux4_1 merge807(
.A0(net1),
.A1(net11),
.A2(net5),
.A3(in44),
.S0(net126),
.S1(net121),
.X(net687)
);

sky130_fd_sc_hd__mux4_4 merge808(
.A0(in0),
.A1(net320),
.A2(net277),
.A3(net462),
.S0(net417),
.S1(net468),
.X(net688)
);

sky130_fd_sc_hd__mux4_4 merge809(
.A0(net230),
.A1(net234),
.A2(net78),
.A3(net114),
.S0(net265),
.S1(net237),
.X(net689)
);

sky130_fd_sc_hd__o221ai_1 merge810(
.A1(net129),
.A2(net147),
.B1(net5),
.B2(net9),
.C1(in58),
.Y(net690)
);

sky130_fd_sc_hd__mux4_4 merge811(
.A0(net81),
.A1(net87),
.A2(net201),
.A3(net203),
.S0(net202),
.S1(net763),
.X(net691)
);

sky130_fd_sc_hd__o221a_1 merge812(
.A1(net121),
.A2(in10),
.B1(in58),
.B2(net123),
.C1(net128),
.X(net692)
);

sky130_fd_sc_hd__mux4_2 merge813(
.A0(net96),
.A1(net142),
.A2(net16),
.A3(net4),
.S0(net19),
.S1(net5),
.X(net693)
);

sky130_fd_sc_hd__mux4_4 merge814(
.A0(net324),
.A1(net311),
.A2(net309),
.A3(in17),
.S0(net200),
.S1(net204),
.X(net694)
);

sky130_fd_sc_hd__mux4_1 merge815(
.A0(net11),
.A1(net16),
.A2(net22),
.A3(net151),
.S0(net140),
.S1(net136),
.X(net695)
);

sky130_fd_sc_hd__mux4_2 merge816(
.A0(net203),
.A1(net199),
.A2(net200),
.A3(in51),
.S0(net233),
.S1(in23),
.X(net696)
);

sky130_fd_sc_hd__mux4_2 merge817(
.A0(net82),
.A1(net317),
.A2(net309),
.A3(net237),
.S0(net220),
.S1(net5),
.X(net697)
);

sky130_fd_sc_hd__mux4_1 merge818(
.A0(net418),
.A1(net450),
.A2(net200),
.A3(net455),
.S0(net453),
.S1(net454),
.X(net698)
);

sky130_fd_sc_hd__mux4_2 merge819(
.A0(out30),
.A1(out53),
.A2(net5),
.A3(net6),
.S0(in10),
.S1(net813),
.X(net699)
);

sky130_fd_sc_hd__mux4_1 merge820(
.A0(net423),
.A1(net424),
.A2(net429),
.A3(net542),
.S0(net535),
.S1(net532),
.X(net700)
);

sky130_fd_sc_hd__mux4_1 merge821(
.A0(in28),
.A1(net80),
.A2(net143),
.A3(net11),
.S0(out30),
.S1(net60),
.X(net701)
);

sky130_fd_sc_hd__mux4_2 merge822(
.A0(net199),
.A1(net309),
.A2(net146),
.A3(net148),
.S0(out52),
.S1(net833),
.X(net702)
);

sky130_fd_sc_hd__o221a_1 merge823(
.A1(net87),
.A2(net205),
.B1(net203),
.B2(net211),
.C1(in21),
.X(net703)
);

sky130_fd_sc_hd__mux4_1 merge824(
.A0(net427),
.A1(net426),
.A2(net432),
.A3(net451),
.S0(net444),
.S1(net449),
.X(net704)
);

sky130_fd_sc_hd__mux4_2 merge825(
.A0(net426),
.A1(net432),
.A2(net428),
.A3(net86),
.S0(net324),
.S1(net430),
.X(net705)
);

sky130_fd_sc_hd__mux4_2 merge826(
.A0(in10),
.A1(net58),
.A2(out30),
.A3(net140),
.S0(net94),
.S1(net25),
.X(net706)
);

sky130_fd_sc_hd__mux4_4 merge827(
.A0(net80),
.A1(net136),
.A2(in12),
.A3(net5),
.S0(net16),
.S1(net740),
.X(net707)
);

sky130_fd_sc_hd__and2b_4 merge828(
.A_N(net456),
.B(net461),
.X(net708)
);

sky130_fd_sc_hd__nand2b_4 merge829(
.A_N(net649),
.B(net691),
.Y(net709)
);

sky130_fd_sc_hd__or2_1 merge830(
.A(net117),
.B(net104),
.X(net710)
);

sky130_fd_sc_hd__dfrbp_1 merge831(
.D(net483),
.RESET_B(net465),
.CLK(clk),
.Q(net712),
.Q_N(net711)
);

sky130_fd_sc_hd__and2_4 merge832(
.A(net300),
.B(net301),
.X(net713)
);

sky130_fd_sc_hd__and2b_2 merge833(
.A_N(net489),
.B(net491),
.X(net714)
);

sky130_fd_sc_hd__nand2_4 merge834(
.A(net269),
.B(net286),
.Y(net715)
);

sky130_fd_sc_hd__and2_2 merge835(
.A(net390),
.B(net391),
.X(net716)
);

sky130_fd_sc_hd__or2_4 merge836(
.A(net630),
.B(net633),
.X(net717)
);

sky130_fd_sc_hd__dfrbp_2 merge837(
.D(net660),
.RESET_B(net677),
.CLK(clk),
.Q(net719),
.Q_N(net718)
);

sky130_fd_sc_hd__nand2b_2 merge838(
.A_N(net590),
.B(net602),
.Y(net720)
);

sky130_fd_sc_hd__dfrtn_1 merge839(
.D(net154),
.RESET_B(net667),
.CLK_N(clk),
.Q(net721)
);

sky130_fd_sc_hd__nand2b_2 merge840(
.A_N(net186),
.B(net189),
.Y(net722)
);

sky130_fd_sc_hd__and2_2 merge841(
.A(net559),
.B(net573),
.X(net723)
);

sky130_fd_sc_hd__nor2_4 merge842(
.A(net515),
.B(net519),
.Y(net724)
);

sky130_fd_sc_hd__dfrtp_1 merge843(
.Q(net46),
.RESET_B(net44),
.CLK(clk)
);

sky130_fd_sc_hd__or2b_1 merge844(
.A(net225),
.B_N(net240),
.X(net726)
);

sky130_fd_sc_hd__nor2b_4 merge845(
.A(net552),
.B_N(net550),
.Y(net727)
);

sky130_fd_sc_hd__dfrtp_2 merge846(
.D(net360),
.RESET_B(net370),
.CLK(clk),
.Q(net728)
);

sky130_fd_sc_hd__dfrtp_4 merge847(
.D(net158),
.RESET_B(net165),
.CLK(clk),
.Q(net729)
);

sky130_fd_sc_hd__or2_2 merge848(
.A(net606),
.B(net607),
.X(net730)
);

sky130_fd_sc_hd__nand2b_1 merge849(
.A_N(net393),
.B(net394),
.Y(net731)
);

sky130_fd_sc_hd__dfsbp_1 merge850(
.D(net659),
.SET_B(net671),
.CLK(clk),
.Q(net733),
.Q_N(net732)
);

sky130_fd_sc_hd__dfsbp_2 merge851(
.D(net650),
.SET_B(net676),
.CLK(clk),
.Q(net735),
.Q_N(net734)
);

sky130_fd_sc_hd__nand2_1 merge852(
.A(net138),
.B(net648),
.Y(net736)
);

sky130_fd_sc_hd__nor2_1 merge853(
.A(net251),
.B(net249),
.Y(net737)
);

sky130_fd_sc_hd__nor2_4 merge854(
.A(net57),
.B(net66),
.Y(net738)
);

sky130_fd_sc_hd__dfstp_1 merge855(
.D(net335),
.SET_B(net339),
.CLK(clk),
.Q(net739)
);

sky130_fd_sc_hd__dfstp_2 merge856(
.D(net10),
.SET_B(net15),
.CLK(clk),
.Q(net740)
);

sky130_fd_sc_hd__dfstp_4 merge857(
.Q(net307),
.SET_B(net306),
.CLK(clk)
);

sky130_fd_sc_hd__nor2b_1 merge858(
.A(net198),
.B_N(net407),
.Y(net741)
);

sky130_fd_sc_hd__dlrbn_1 merge859(
.D(net702),
.RESET_B(net644),
.GATE_N(clk),
.Q(net743),
.Q_N(net742)
);

sky130_fd_sc_hd__and2b_2 merge860(
.A_N(net197),
.B(net194),
.X(net744)
);

sky130_fd_sc_hd__dlrbn_2 merge861(
.D(net694),
.RESET_B(net683),
.GATE_N(clk),
.Q(net746),
.Q_N(net745)
);

sky130_fd_sc_hd__and2b_1 merge862(
.A_N(net287),
.B(net713),
.X(net747)
);

sky130_fd_sc_hd__dlrbp_1 merge863(
.D(net678),
.RESET_B(net696),
.GATE(clk),
.Q(net749),
.Q_N(net748)
);

sky130_fd_sc_hd__or2_1 merge864(
.A(net618),
.B(net642),
.X(net750)
);

sky130_fd_sc_hd__dlrbp_2 merge865(
.D(net708),
.RESET_B(net703),
.GATE(clk),
.Q(net752),
.Q_N(net751)
);

sky130_fd_sc_hd__nor2b_4 merge866(
.A(net574),
.B_N(net578),
.Y(net753)
);

sky130_fd_sc_hd__and2b_1 merge867(
.A_N(net525),
.B(net640),
.X(net754)
);

sky130_fd_sc_hd__and2b_4 merge868(
.A_N(net400),
.B(net415),
.X(net755)
);

sky130_fd_sc_hd__or2b_4 merge869(
.A(net608),
.B_N(net639),
.X(net756)
);

sky130_fd_sc_hd__and2b_4 merge870(
.A_N(net501),
.B(net527),
.X(net757)
);

sky130_fd_sc_hd__dlrtn_1 merge871(
.D(net604),
.RESET_B(net720),
.GATE_N(clk),
.Q(net758)
);

sky130_fd_sc_hd__dlrtn_2 merge872(
.D(net647),
.RESET_B(net684),
.GATE_N(clk),
.Q(net759)
);

sky130_fd_sc_hd__dlrtn_4 merge873(
.D(net657),
.RESET_B(net675),
.GATE_N(clk),
.Q(net760)
);

sky130_fd_sc_hd__dlrtp_1 merge874(
.D(net680),
.RESET_B(net723),
.GATE(clk),
.Q(net761)
);

sky130_fd_sc_hd__or2_1 merge875(
.A(net619),
.B(net506),
.X(net762)
);

sky130_fd_sc_hd__dlrtp_2 merge876(
.D(net692),
.RESET_B(net84),
.GATE(clk),
.Q(net763)
);

sky130_fd_sc_hd__nand2b_1 merge877(
.A_N(net399),
.B(net523),
.Y(net764)
);

sky130_fd_sc_hd__dlrtp_4 merge878(
.D(net710),
.RESET_B(net709),
.GATE(clk),
.Q(net765)
);

sky130_fd_sc_hd__nor2_4 merge879(
.A(net520),
.B(net625),
.Y(net766)
);

sky130_fd_sc_hd__edfxbp_1 merge880(
.D(net193),
.DE(net302),
.CLK(clk),
.Q(out49),
.Q_N(net767)
);

sky130_fd_sc_hd__edfxtp_1 merge881(
.D(net652),
.DE(net655),
.CLK(clk),
.Q(net768)
);

sky130_fd_sc_hd__sdlclkp_1 merge882(
.GATE(net166),
.SCE(net687),
.CLK(clk),
.GCLK(net769)
);

sky130_fd_sc_hd__sdlclkp_2 merge883(
.GATE(net611),
.SCE(net624),
.CLK(clk),
.GCLK(net770)
);

sky130_fd_sc_hd__sdlclkp_4 merge884(
.GATE(net681),
.SCE(net695),
.CLK(clk),
.GCLK(net771)
);

sky130_fd_sc_hd__dfrbp_1 merge885(
.D(net658),
.RESET_B(net727),
.CLK(clk),
.Q(net773),
.Q_N(net772)
);

sky130_fd_sc_hd__dfrbp_2 merge886(
.D(net755),
.RESET_B(net289),
.CLK(clk),
.Q(out12),
.Q_N(net774)
);

sky130_fd_sc_hd__dfrtn_1 merge887(
.D(net651),
.RESET_B(net679),
.CLK_N(clk),
.Q(net775)
);

sky130_fd_sc_hd__dfrtp_1 merge888(
.D(net697),
.RESET_B(net682),
.CLK(clk),
.Q(net776)
);

sky130_fd_sc_hd__dfrtp_2 merge889(
.D(net716),
.RESET_B(net701),
.CLK(clk),
.Q(net777)
);

sky130_fd_sc_hd__dfrtp_4 merge890(
.D(net715),
.RESET_B(net668),
.CLK(clk),
.Q(net778)
);

sky130_fd_sc_hd__dfsbp_1 merge891(
.D(net177),
.SET_B(net744),
.CLK(clk),
.Q(net779),
.Q_N(out57)
);

sky130_fd_sc_hd__dfsbp_2 merge892(
.D(net511),
.SET_B(net514),
.CLK(clk),
.Q(net781),
.Q_N(net780)
);

sky130_fd_sc_hd__nand2_4 merge893(
.A(net613),
.B(net623),
.Y(net782)
);

sky130_fd_sc_hd__nor2_1 merge894(
.A(net622),
.B(net615),
.Y(net783)
);

sky130_fd_sc_hd__dfstp_1 merge895(
.D(net665),
.SET_B(net741),
.CLK(clk),
.Q(net784)
);

sky130_fd_sc_hd__dfstp_2 merge896(
.D(net621),
.SET_B(net663),
.CLK(clk),
.Q(net785)
);

sky130_fd_sc_hd__dfstp_4 merge897(
.D(net653),
.SET_B(net689),
.CLK(clk),
.Q(net786)
);

sky130_fd_sc_hd__dlrbn_1 merge898(
.D(net690),
.RESET_B(net722),
.GATE_N(clk),
.Q(net788),
.Q_N(net787)
);

sky130_fd_sc_hd__dlrbn_2 merge899(
.D(net693),
.RESET_B(net706),
.GATE_N(clk),
.Q(net790),
.Q_N(net789)
);

sky130_fd_sc_hd__dlrbp_1 merge900(
.D(net700),
.RESET_B(net605),
.GATE(clk),
.Q(net792),
.Q_N(net791)
);

sky130_fd_sc_hd__dlrbp_2 merge901(
.D(net279),
.RESET_B(net699),
.GATE(clk),
.Q(net794),
.Q_N(net793)
);

sky130_fd_sc_hd__dlrtn_1 merge902(
.D(net753),
.RESET_B(net603),
.GATE_N(clk),
.Q(net795)
);

sky130_fd_sc_hd__dlrtn_2 merge903(
.D(net717),
.RESET_B(net766),
.GATE_N(clk),
.Q(net796)
);

sky130_fd_sc_hd__dlrtn_4 merge904(
.D(net349),
.RESET_B(net344),
.GATE_N(clk),
.Q(net797)
);

sky130_fd_sc_hd__dlrtp_1 merge905(
.D(net730),
.RESET_B(net662),
.GATE(clk),
.Q(net798)
);

sky130_fd_sc_hd__dlrtp_2 merge906(
.D(net466),
.RESET_B(net591),
.GATE(clk),
.Q(net799)
);

sky130_fd_sc_hd__dlrtp_4 merge907(
.D(net477),
.RESET_B(net688),
.GATE(clk),
.Q(net800)
);

sky130_fd_sc_hd__edfxbp_1 merge908(
.D(net268),
.DE(net698),
.CLK(clk),
.Q(net802),
.Q_N(net801)
);

sky130_fd_sc_hd__edfxtp_1 merge909(
.D(net750),
.DE(net754),
.CLK(clk),
.Q(net803)
);

sky130_fd_sc_hd__sdlclkp_1 merge910(
.GATE(net757),
.SCE(net670),
.CLK(clk),
.GCLK(out15)
);

sky130_fd_sc_hd__sdlclkp_2 merge911(
.GATE(net666),
.SCE(net664),
.CLK(clk),
.GCLK(net804)
);

sky130_fd_sc_hd__sdlclkp_4 merge912(
.GATE(net686),
.SCE(net196),
.CLK(clk),
.GCLK(net805)
);

sky130_fd_sc_hd__dfrbp_1 merge913(
.D(net704),
.RESET_B(net705),
.CLK(clk),
.Q(net807),
.Q_N(net806)
);

sky130_fd_sc_hd__dfrbp_2 merge914(
.D(net397),
.RESET_B(net672),
.CLK(clk),
.Q(net809),
.Q_N(net808)
);

sky130_fd_sc_hd__dfrtn_1 merge915(
.D(net707),
.RESET_B(net738),
.CLK_N(clk),
.Q(net810)
);

sky130_fd_sc_hd__dfrtp_1 merge916(
.D(net510),
.RESET_B(net502),
.CLK(clk),
.Q(net811)
);

sky130_fd_sc_hd__dfrtp_2 merge917(
.D(net726),
.RESET_B(net747),
.CLK(clk),
.Q(net812)
);

sky130_fd_sc_hd__dfrtp_4 merge918(
.D(net63),
.RESET_B(net674),
.CLK(clk),
.Q(net813)
);

sky130_fd_sc_hd__dfsbp_1 merge919(
.D(net714),
.SET_B(net656),
.CLK(clk),
.Q(out8),
.Q_N(net814)
);

sky130_fd_sc_hd__dfsbp_2 merge920(
.D(net764),
.SET_B(net731),
.CLK(clk),
.Q(net815),
.Q_N(out14)
);

sky130_fd_sc_hd__dfstp_1 merge921(
.D(net685),
.SET_B(net724),
.CLK(clk),
.Q(net816)
);

sky130_fd_sc_hd__dfstp_2 merge922(
.D(net582),
.SET_B(net673),
.CLK(clk),
.Q(net817)
);

sky130_fd_sc_hd__dfstp_4 merge923(
.D(net325),
.SET_B(net384),
.CLK(clk),
.Q(net818)
);

sky130_fd_sc_hd__dlrbn_1 merge924(
.D(net736),
.RESET_B(net737),
.GATE_N(clk),
.Q(net820),
.Q_N(net819)
);

sky130_fd_sc_hd__dlrbn_2 merge925(
.D(net783),
.RESET_B(net782),
.GATE_N(clk),
.Q(net822),
.Q_N(net821)
);

sky130_fd_sc_hd__dlrbp_1 merge926(
.D(net398),
.RESET_B(net499),
.GATE(clk),
.Q(net823),
.Q_N(out9)
);

sky130_fd_sc_hd__dlrbp_2 merge927(
.D(net518),
.RESET_B(net756),
.GATE(clk),
.Q(net825),
.Q_N(net824)
);

sky130_fd_sc_hd__dlrtn_1 merge928(
.D(net517),
.RESET_B(net762),
.GATE_N(clk),
.Q(out11)
);

sky130_fd_sc_hd__dlrtn_2 merge929(
.D(net414),
.RESET_B(net405),
.GATE_N(clk),
.Q(out25)
);

sky130_fd_sc_hd__dfxbp_1 s930(
.D(net40),
.CLK(clk),
.Q(net827),
.Q_N(net826)
);

sky130_fd_sc_hd__dfxbp_2 s931(
.D(net68),
.CLK(clk),
.Q(out31),
.Q_N(net828)
);

sky130_fd_sc_hd__dfxtp_1 s932(
.D(net116),
.CLK(clk),
.Q(net829)
);

sky130_fd_sc_hd__dfxtp_2 s933(
.D(net134),
.CLK(clk),
.Q(net830)
);

sky130_fd_sc_hd__dfxtp_4 s934(
.D(net137),
.CLK(clk),
.Q(net831)
);

sky130_fd_sc_hd__dlclkp_1 s935(
.GATE(net155),
.CLK(clk),
.GCLK(net832)
);

sky130_fd_sc_hd__dlclkp_2 s936(
.GATE(net156),
.CLK(clk),
.GCLK(out4)
);

sky130_fd_sc_hd__dlclkp_4 s937(
.GATE(net188),
.CLK(clk),
.GCLK(out54)
);

sky130_fd_sc_hd__dlxbn_1 s938(
.D(net219),
.GATE_N(clk),
.Q(net834),
.Q_N(net833)
);

sky130_fd_sc_hd__dlxbn_2 s939(
.D(net222),
.GATE_N(clk),
.Q(out0),
.Q_N(net835)
);

sky130_fd_sc_hd__dlxbp_1 s940(
.D(net243),
.GATE(clk),
.Q(net837),
.Q_N(net836)
);

sky130_fd_sc_hd__dlxtn_1 s941(
.D(net250),
.GATE_N(clk),
.Q(net838)
);

sky130_fd_sc_hd__dlxtn_2 s942(
.D(net253),
.GATE_N(clk),
.Q(net839)
);

sky130_fd_sc_hd__dlxtn_4 s943(
.D(net282),
.GATE_N(clk),
.Q(net840)
);

sky130_fd_sc_hd__dlxtp_1 s944(
.D(net285),
.GATE(clk),
.Q(net841)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s945(
.D(net288),
.SLEEP_B(clk),
.Q(net842)
);

sky130_fd_sc_hd__dfxbp_1 s946(
.D(net295),
.CLK(clk),
.Q(net844),
.Q_N(net843)
);

sky130_fd_sc_hd__dfxbp_2 s947(
.D(net299),
.CLK(clk),
.Q(net846),
.Q_N(net845)
);

sky130_fd_sc_hd__dfxtp_1 s948(
.D(net305),
.CLK(clk),
.Q(out29)
);

sky130_fd_sc_hd__dfxtp_2 s949(
.D(net323),
.CLK(clk),
.Q(out38)
);

sky130_fd_sc_hd__dfxtp_4 s950(
.D(net327),
.CLK(clk),
.Q(net847)
);

sky130_fd_sc_hd__dlclkp_1 s951(
.GATE(net328),
.CLK(clk),
.GCLK(net848)
);

sky130_fd_sc_hd__dlclkp_2 s952(
.GATE(net340),
.CLK(clk),
.GCLK(net849)
);

sky130_fd_sc_hd__dlclkp_4 s953(
.GATE(net343),
.CLK(clk),
.GCLK(net850)
);

sky130_fd_sc_hd__dlxbn_1 s954(
.D(net345),
.GATE_N(clk),
.Q(net852),
.Q_N(net851)
);

sky130_fd_sc_hd__dlxbn_2 s955(
.D(net346),
.GATE_N(clk),
.Q(net854),
.Q_N(net853)
);

sky130_fd_sc_hd__dlxbp_1 s956(
.D(net348),
.GATE(clk),
.Q(net856),
.Q_N(net855)
);

sky130_fd_sc_hd__dlxtn_1 s957(
.D(net368),
.GATE_N(clk),
.Q(net857)
);

sky130_fd_sc_hd__dlxtn_2 s958(
.D(net369),
.GATE_N(clk),
.Q(out3)
);

sky130_fd_sc_hd__dlxtn_4 s959(
.D(net406),
.GATE_N(clk),
.Q(net858)
);

sky130_fd_sc_hd__dlxtp_1 s960(
.D(net408),
.GATE(clk),
.Q(net859)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s961(
.D(net412),
.SLEEP_B(clk),
.Q(net860)
);

sky130_fd_sc_hd__dfxbp_1 s962(
.D(net435),
.CLK(clk),
.Q(net862),
.Q_N(net861)
);

sky130_fd_sc_hd__dfxbp_2 s963(
.D(net472),
.CLK(clk),
.Q(net864),
.Q_N(net863)
);

sky130_fd_sc_hd__dfxtp_1 s964(
.D(net474),
.CLK(clk),
.Q(net865)
);

sky130_fd_sc_hd__dfxtp_2 s965(
.D(net475),
.CLK(clk),
.Q(net866)
);

sky130_fd_sc_hd__dfxtp_4 s966(
.D(net482),
.CLK(clk),
.Q(net867)
);

sky130_fd_sc_hd__dlclkp_1 s967(
.GATE(net486),
.CLK(clk),
.GCLK(net868)
);

sky130_fd_sc_hd__dlclkp_2 s968(
.GATE(net490),
.CLK(clk),
.GCLK(net869)
);

sky130_fd_sc_hd__dlclkp_4 s969(
.GATE(net493),
.CLK(clk),
.GCLK(out17)
);

sky130_fd_sc_hd__dlxbn_1 s970(
.D(net505),
.GATE_N(clk),
.Q(net871),
.Q_N(net870)
);

sky130_fd_sc_hd__dlxbn_2 s971(
.D(net507),
.GATE_N(clk),
.Q(net873),
.Q_N(net872)
);

sky130_fd_sc_hd__dlxbp_1 s972(
.D(net512),
.GATE(clk),
.Q(net875),
.Q_N(net874)
);

sky130_fd_sc_hd__dlxtn_1 s973(
.D(net524),
.GATE_N(clk),
.Q(out20)
);

sky130_fd_sc_hd__dlxtn_2 s974(
.D(net526),
.GATE_N(clk),
.Q(net876)
);

sky130_fd_sc_hd__dlxtn_4 s975(
.D(net529),
.GATE_N(clk),
.Q(net877)
);

sky130_fd_sc_hd__dlxtp_1 s976(
.D(net531),
.GATE(clk),
.Q(net878)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s977(
.D(net544),
.SLEEP_B(clk),
.Q(net879)
);

sky130_fd_sc_hd__dfxbp_1 s978(
.D(net563),
.CLK(clk),
.Q(net881),
.Q_N(net880)
);

sky130_fd_sc_hd__dfxbp_2 s979(
.D(net571),
.CLK(clk),
.Q(net883),
.Q_N(net882)
);

sky130_fd_sc_hd__dfxtp_1 s980(
.D(net583),
.CLK(clk),
.Q(net884)
);

sky130_fd_sc_hd__dfxtp_2 s981(
.D(net592),
.CLK(clk),
.Q(net885)
);

sky130_fd_sc_hd__dfxtp_4 s982(
.D(net600),
.CLK(clk),
.Q(net886)
);

sky130_fd_sc_hd__dlclkp_1 s983(
.GATE(net609),
.CLK(clk),
.GCLK(net887)
);

sky130_fd_sc_hd__dlclkp_2 s984(
.GATE(net610),
.CLK(clk),
.GCLK(net888)
);

sky130_fd_sc_hd__dlclkp_4 s985(
.GATE(net614),
.CLK(clk),
.GCLK(net889)
);

sky130_fd_sc_hd__dlxbn_1 s986(
.D(net620),
.GATE_N(clk),
.Q(net891),
.Q_N(net890)
);

sky130_fd_sc_hd__dlxbn_2 s987(
.D(net626),
.GATE_N(clk),
.Q(net893),
.Q_N(net892)
);

sky130_fd_sc_hd__dlxbp_1 s988(
.D(net627),
.GATE(clk),
.Q(net895),
.Q_N(net894)
);

sky130_fd_sc_hd__dlxtn_1 s989(
.D(net635),
.GATE_N(clk),
.Q(net896)
);

sky130_fd_sc_hd__dlxtn_2 s990(
.D(net637),
.GATE_N(clk),
.Q(net897)
);


endmodule
