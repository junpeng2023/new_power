module netlist_4 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51
);


wire net664;
wire net659;
wire net656;
wire net652;
wire net651;
wire net645;
wire net641;
wire net637;
wire net632;
wire out18;
wire net631;
wire net629;
wire net628;
wire net627;
wire net626;
wire net624;
wire net623;
wire net620;
wire net619;
wire net615;
wire out17;
wire net614;
wire net613;
wire net612;
wire net638;
wire net610;
wire net608;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire out1;
wire out7;
wire net596;
wire net595;
wire net592;
wire net588;
wire net587;
wire net583;
wire net582;
wire net584;
wire net581;
wire net579;
wire net577;
wire net576;
wire net569;
wire net567;
wire net566;
wire net565;
wire net562;
wire net559;
wire net556;
wire net647;
wire net555;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire net550;
wire net544;
wire net539;
wire net534;
wire net532;
wire net530;
wire net617;
wire net537;
wire net528;
wire net525;
wire net523;
wire net520;
wire net519;
wire net516;
wire net514;
wire net508;
wire net504;
wire net503;
wire net499;
wire clk;
wire net496;
wire net495;
wire net494;
wire net493;
wire net492;
wire net491;
wire net490;
wire net489;
wire net487;
wire net486;
wire net478;
wire net474;
wire net473;
wire net472;
wire net468;
wire net540;
wire net465;
wire net462;
wire net469;
wire net461;
wire net546;
wire net460;
wire net454;
wire net453;
wire net648;
wire net452;
wire net449;
wire net448;
wire net498;
wire net446;
wire net444;
wire net442;
wire out15;
wire net441;
wire net609;
wire net440;
wire net439;
wire net438;
wire net433;
wire net432;
wire net431;
wire net430;
wire net618;
wire net429;
wire net428;
wire net427;
wire net570;
wire out2;
wire out49;
wire out48;
wire out13;
wire net426;
wire net425;
wire net423;
wire net531;
wire net421;
wire net420;
wire out38;
wire net450;
wire net418;
wire out33;
wire net416;
wire net415;
wire net414;
wire net413;
wire net412;
wire net411;
wire net410;
wire net409;
wire out26;
wire net408;
wire net407;
wire net662;
wire net405;
wire out37;
wire net607;
wire net526;
wire net404;
wire net403;
wire net663;
wire net402;
wire net572;
wire net401;
wire out46;
wire net399;
wire net406;
wire out19;
wire net398;
wire net476;
wire net396;
wire out3;
wire net395;
wire net391;
wire net557;
wire net527;
wire net488;
wire net390;
wire net646;
wire net389;
wire net513;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net380;
wire net379;
wire net616;
wire net378;
wire net377;
wire net376;
wire net580;
wire net375;
wire net625;
wire net598;
wire net374;
wire net373;
wire net372;
wire net371;
wire net370;
wire net368;
wire net367;
wire net366;
wire net365;
wire net364;
wire net363;
wire net360;
wire net397;
wire net357;
wire net356;
wire net355;
wire out25;
wire net521;
wire net353;
wire net590;
wire net507;
wire net351;
wire net350;
wire net547;
wire net511;
wire net343;
wire net348;
wire net341;
wire net340;
wire net339;
wire net337;
wire net336;
wire net538;
wire net334;
wire net333;
wire net332;
wire net331;
wire out32;
wire net330;
wire net517;
wire net328;
wire net327;
wire net325;
wire net324;
wire net299;
wire net143;
wire net322;
wire net505;
wire net312;
wire net319;
wire net318;
wire out43;
wire net342;
wire net17;
wire out44;
wire net636;
wire in37;
wire net159;
wire net311;
wire out14;
wire net309;
wire net417;
wire out8;
wire net302;
wire net298;
wire net296;
wire in24;
wire net295;
wire net358;
wire net127;
wire net294;
wire in49;
wire net147;
wire net180;
wire net310;
wire net293;
wire net305;
wire out39;
wire in4;
wire net292;
wire net500;
wire net445;
wire out22;
wire net291;
wire net665;
wire net422;
wire net289;
wire net482;
wire in25;
wire net288;
wire net589;
wire net424;
wire net278;
wire net276;
wire net274;
wire net643;
wire net273;
wire out10;
wire in39;
wire net272;
wire net114;
wire net270;
wire in17;
wire net267;
wire net644;
wire net266;
wire net463;
wire net297;
wire net475;
wire out27;
wire net102;
wire net151;
wire net264;
wire net657;
wire net591;
wire net262;
wire net217;
wire net261;
wire net257;
wire net117;
wire net62;
wire net254;
wire net203;
wire net253;
wire net252;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire net111;
wire net242;
wire net661;
wire net241;
wire net573;
wire net240;
wire out42;
wire net238;
wire net142;
wire net183;
wire net234;
wire net232;
wire out12;
wire net226;
wire net244;
wire net568;
wire net223;
wire net524;
wire net382;
wire net259;
wire net335;
wire net222;
wire net219;
wire net578;
wire net210;
wire net213;
wire net208;
wire out16;
wire net188;
wire net207;
wire net649;
wire net205;
wire net202;
wire net130;
wire net201;
wire net384;
wire net224;
wire net122;
wire net197;
wire net193;
wire net192;
wire net190;
wire in35;
wire out24;
wire in20;
wire net189;
wire net246;
wire net186;
wire net164;
wire out0;
wire net126;
wire net284;
wire net655;
wire net563;
wire net549;
wire net182;
wire net133;
wire net175;
wire net173;
wire net195;
wire net479;
wire net8;
wire net172;
wire net622;
wire net518;
wire net170;
wire net381;
wire net218;
wire net169;
wire net344;
wire net168;
wire net286;
wire net167;
wire net58;
wire net221;
wire net166;
wire net269;
wire net165;
wire net660;
wire net359;
wire out28;
wire net575;
wire net434;
wire net200;
wire net162;
wire net497;
wire out45;
wire net161;
wire net316;
wire out31;
wire net285;
wire net160;
wire net158;
wire net152;
wire net150;
wire net149;
wire net148;
wire net178;
wire net239;
wire net144;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net561;
wire out29;
wire net139;
wire net5;
wire out41;
wire net456;
wire net135;
wire net157;
wire net177;
wire out51;
wire net134;
wire in12;
wire net271;
wire net103;
wire net124;
wire net255;
wire net548;
wire net481;
wire net383;
wire net120;
wire net100;
wire net455;
wire net129;
wire net392;
wire net113;
wire net204;
wire net110;
wire net109;
wire net642;
wire net268;
wire in7;
wire net82;
wire net123;
wire net282;
wire net71;
wire net229;
wire net326;
wire net108;
wire net107;
wire net104;
wire net99;
wire net96;
wire net225;
wire net250;
wire net466;
wire net118;
wire net94;
wire net90;
wire net74;
wire net277;
wire net639;
wire net88;
wire net81;
wire net230;
wire net156;
wire net361;
wire net115;
wire net209;
wire net258;
wire out40;
wire in18;
wire net34;
wire net79;
wire net75;
wire net306;
wire net231;
wire net349;
wire net329;
wire net212;
wire net653;
wire net485;
wire net78;
wire in5;
wire net77;
wire net236;
wire net76;
wire net354;
wire in38;
wire net198;
wire net467;
wire net101;
wire out20;
wire net9;
wire net136;
wire net571;
wire net31;
wire net73;
wire net199;
wire out21;
wire net60;
wire net179;
wire net564;
wire net443;
wire net154;
wire net345;
wire net84;
wire in46;
wire net85;
wire net72;
wire net116;
wire net69;
wire net128;
wire net67;
wire in31;
wire net65;
wire net447;
wire net98;
wire net522;
wire net459;
wire net436;
wire out9;
wire net260;
wire net541;
wire net501;
wire net323;
wire net15;
wire net64;
wire net63;
wire net61;
wire net512;
wire out34;
wire net237;
wire net59;
wire net248;
wire net275;
wire net119;
wire net477;
wire net400;
wire in10;
wire net57;
wire net228;
wire net39;
wire net630;
wire net56;
wire net55;
wire net214;
wire net53;
wire net97;
wire in48;
wire net196;
wire net52;
wire net640;
wire net369;
wire net50;
wire net597;
wire net155;
wire net338;
wire net46;
wire net599;
wire net112;
wire net650;
wire net185;
wire net585;
wire net560;
wire net45;
wire net502;
wire net235;
wire net49;
wire net594;
wire net215;
wire net484;
wire net184;
wire out36;
wire in8;
wire net346;
wire net43;
wire net435;
wire net18;
wire net121;
wire net304;
wire net40;
wire net437;
wire in36;
wire out30;
wire net558;
wire in1;
wire net13;
wire net265;
wire net457;
wire out4;
wire net91;
wire net42;
wire net536;
wire net37;
wire net27;
wire net54;
wire net281;
wire net36;
wire net21;
wire net35;
wire net187;
wire in13;
wire net621;
wire net586;
wire net533;
wire net32;
wire net419;
wire net125;
wire net458;
wire net19;
wire net347;
wire in15;
wire net20;
wire in19;
wire net70;
wire net48;
wire net28;
wire net92;
wire net25;
wire net30;
wire net29;
wire in0;
wire net24;
wire net263;
wire out50;
wire net6;
wire net315;
wire net22;
wire net464;
wire net3;
wire net176;
wire out23;
wire out47;
wire net290;
wire net227;
wire net470;
wire net44;
wire net471;
wire in33;
wire net33;
wire net233;
wire net535;
wire net320;
wire net301;
wire net26;
wire net483;
wire net16;
wire in28;
wire net41;
wire out11;
wire net206;
wire net138;
wire net211;
wire in6;
wire net0;
wire net132;
wire net106;
wire net303;
wire in34;
wire net593;
wire in45;
wire net163;
wire net393;
wire net4;
wire in42;
wire net321;
wire net256;
wire net87;
wire net509;
wire net506;
wire net181;
wire net451;
wire net7;
wire net145;
wire net574;
wire net23;
wire net216;
wire out5;
wire net14;
wire net2;
wire in44;
wire net601;
wire out35;
wire in32;
wire in50;
wire net47;
wire net12;
wire in27;
wire in9;
wire net654;
wire net611;
wire net515;
wire net362;
wire in16;
wire net191;
wire net89;
wire in41;
wire in26;
wire net543;
wire net220;
wire net171;
wire in43;
wire net174;
wire in22;
wire net308;
wire out6;
wire net600;
wire net510;
wire net68;
wire in14;
wire net529;
wire in21;
wire net480;
wire net86;
wire net317;
wire in51;
wire net93;
wire net280;
wire in47;
wire net137;
wire in2;
wire net131;
wire net658;
wire net105;
wire in11;
wire net38;
wire net51;
wire net153;
wire net95;
wire net300;
wire in30;
wire net146;
wire net279;
wire in23;
wire net394;
wire in3;
wire net314;
wire net251;
wire net11;
wire net352;
wire net307;
wire net633;
wire net194;
wire net542;
wire net80;
wire in29;
wire net313;
wire net1;
sky130_fd_sc_hd__a21boi_0 c52(
.A1(in30),
.A2(in50),
.B1_N(in51),
.Y(net0)
);

sky130_fd_sc_hd__a21oi_2 c53(
.A1(in49),
.A2(in24),
.B1(in51),
.Y(net1)
);

sky130_fd_sc_hd__o41a_2 c54(
.A1(net0),
.A2(in44),
.A3(net1),
.A4(in43),
.B1(in51),
.X(net2)
);

sky130_fd_sc_hd__a21o_1 c55(
.A1(in46),
.A2(in42),
.B1(in47),
.X(net3)
);

sky130_fd_sc_hd__o41a_1 c56(
.A1(in36),
.A2(net3),
.A3(in45),
.A4(in38),
.B1(in51),
.X(net4)
);

sky130_fd_sc_hd__o21ai_0 c57(
.A1(in47),
.A2(in50),
.B1(net2),
.Y(net5)
);

sky130_fd_sc_hd__o31ai_2 c58(
.A1(net4),
.A2(in21),
.A3(in30),
.B1(in51),
.Y(net6)
);

sky130_fd_sc_hd__a21o_1 c59(
.A1(in42),
.A2(in45),
.B1(net6),
.X(net7)
);

sky130_fd_sc_hd__o21ai_0 c60(
.A1(net5),
.A2(in40),
.B1(in21),
.Y(net8)
);

sky130_fd_sc_hd__o21ba_4 c61(
.A1(in21),
.A2(net7),
.B1_N(net4),
.X(net9)
);

sky130_fd_sc_hd__o21ai_0 c62(
.A1(net8),
.A2(net9),
.B1(in2),
.Y(net10)
);

sky130_fd_sc_hd__or2_2 c63(
.A(in38),
.B(net12),
.X(net11)
);

sky130_fd_sc_hd__nor2b_1 c64(
.A(in46),
.B_N(net5),
.Y(out11)
);

sky130_fd_sc_hd__and2_0 c65(
.A(in15),
.B(in7),
.X(net12)
);

sky130_fd_sc_hd__or2b_2 c66(
.A(net6),
.B_N(in46),
.X(net13)
);

sky130_fd_sc_hd__or2_4 c67(
.A(in16),
.B(net5),
.X(net14)
);

sky130_fd_sc_hd__nor2_4 c68(
.A(net13),
.B(net1),
.Y(net15)
);

sky130_fd_sc_hd__and2_4 c69(
.A(in2),
.B(out11),
.X(net16)
);

sky130_fd_sc_hd__and2_1 c70(
.A(out11),
.B(net11),
.X(net17)
);

sky130_fd_sc_hd__nor2_4 c71(
.A(net11),
.B(in19),
.Y(net18)
);

sky130_fd_sc_hd__a21boi_2 c72(
.A1(in24),
.A2(net18),
.B1_N(out11),
.Y(net19)
);

sky130_fd_sc_hd__and2_1 c73(
.A(net19),
.B(net16),
.X(net20)
);

sky130_fd_sc_hd__o21bai_4 c74(
.A1(net14),
.A2(net17),
.B1_N(net19),
.Y(net21)
);

sky130_fd_sc_hd__or2b_1 c75(
.A(net20),
.B_N(net21),
.X(net22)
);

sky130_fd_sc_hd__and2_1 c76(
.A(net18),
.B(net19),
.X(net23)
);

sky130_fd_sc_hd__mux2_1 c77(
.A0(net13),
.A1(in39),
.S(in38),
.X(net24)
);

sky130_fd_sc_hd__and2b_2 c78(
.A_N(net16),
.B(net19),
.X(net25)
);

sky130_fd_sc_hd__nor2_1 c79(
.A(net25),
.B(net15),
.Y(net26)
);

sky130_fd_sc_hd__o31ai_1 c80(
.A1(in44),
.A2(net22),
.A3(net26),
.B1(net25),
.Y(net27)
);

sky130_fd_sc_hd__o31ai_1 c81(
.A1(net21),
.A2(net27),
.A3(net23),
.B1(in2),
.Y(out6)
);

sky130_fd_sc_hd__o21ai_4 c82(
.A1(net26),
.A2(net25),
.B1(net20),
.Y(net28)
);

sky130_fd_sc_hd__o31ai_2 c83(
.A1(net22),
.A2(net27),
.A3(net21),
.B1(in51),
.Y(net29)
);

sky130_fd_sc_hd__buf_8 c84(
.A(net25),
.X(net30)
);

sky130_fd_sc_hd__clkinv_2 c85(
.A(in39),
.Y(net31)
);

sky130_fd_sc_hd__buf_6 c86(
.A(net7),
.X(net32)
);

sky130_fd_sc_hd__or2b_1 c87(
.A(net30),
.B_N(net32),
.X(net33)
);

sky130_fd_sc_hd__nand2_4 c88(
.A(in49),
.B(net12),
.Y(net34)
);

sky130_fd_sc_hd__or2_2 c89(
.A(net30),
.B(net11),
.X(net35)
);

sky130_fd_sc_hd__nor2_4 c90(
.A(net9),
.B(net3),
.Y(net36)
);

sky130_fd_sc_hd__nand2_2 c91(
.A(net35),
.B(net30),
.Y(net37)
);

sky130_fd_sc_hd__and2_4 c92(
.A(net34),
.B(net36),
.X(net38)
);

sky130_fd_sc_hd__and2_4 c93(
.A(net35),
.B(net34),
.X(net39)
);

sky130_fd_sc_hd__o21bai_4 c94(
.A1(net3),
.A2(net36),
.B1_N(net12),
.Y(net40)
);

sky130_fd_sc_hd__nand2b_4 c95(
.A_N(net40),
.B(net36),
.Y(net41)
);

sky130_fd_sc_hd__nor2_2 c96(
.A(net36),
.B(net38),
.Y(net42)
);

sky130_fd_sc_hd__or2_4 c97(
.A(net37),
.B(net39),
.X(net43)
);

sky130_fd_sc_hd__nor2_1 c98(
.A(net43),
.B(net15),
.Y(net44)
);

sky130_fd_sc_hd__nand2b_4 c99(
.A_N(net44),
.B(net14),
.Y(net45)
);

sky130_fd_sc_hd__o21bai_4 c100(
.A1(net45),
.A2(net44),
.B1_N(net35),
.Y(net46)
);

sky130_fd_sc_hd__a21boi_2 c101(
.A1(in22),
.A2(net43),
.B1_N(net39),
.Y(net47)
);

sky130_fd_sc_hd__and2_4 c102(
.A(net47),
.B(net32),
.X(net48)
);

sky130_fd_sc_hd__a21bo_1 c103(
.A1(net41),
.A2(net47),
.B1_N(net46),
.X(net49)
);

sky130_fd_sc_hd__mux4_1 c104(
.A0(net32),
.A1(net19),
.A2(net7),
.A3(net48),
.S0(net47),
.S1(in51),
.X(net50)
);

sky130_fd_sc_hd__nand2_4 c105(
.A(in42),
.B(net48),
.Y(net51)
);

sky130_fd_sc_hd__nand2b_1 c106(
.A_N(net4),
.B(net5),
.Y(net52)
);

sky130_fd_sc_hd__o21ai_0 c107(
.A1(net5),
.A2(net48),
.B1(in51),
.Y(out34)
);

sky130_fd_sc_hd__or2_1 c108(
.A(net51),
.B(net11),
.X(net53)
);

sky130_fd_sc_hd__nor2b_2 c109(
.A(out34),
.B_N(net53),
.Y(net54)
);

sky130_fd_sc_hd__or2_2 c110(
.A(net53),
.B(net0),
.X(net55)
);

sky130_fd_sc_hd__dfrbp_1 c111(
.D(net55),
.RESET_B(net47),
.CLK(clk),
.Q(net57),
.Q_N(net56)
);

sky130_fd_sc_hd__or2_1 c112(
.A(in47),
.B(net53),
.X(net58)
);

sky130_fd_sc_hd__nand2_1 c113(
.A(net0),
.B(net42),
.Y(net59)
);

sky130_fd_sc_hd__dfrbp_2 c114(
.D(net54),
.RESET_B(net0),
.CLK(clk),
.Q(net61),
.Q_N(net60)
);

sky130_fd_sc_hd__dfrtn_1 c115(
.D(net54),
.RESET_B(net58),
.CLK_N(clk),
.Q(net62)
);

sky130_fd_sc_hd__nor2_1 c116(
.A(in45),
.B(net56),
.Y(net63)
);

sky130_fd_sc_hd__nor2_4 c117(
.A(net59),
.B(net63),
.Y(net64)
);

sky130_fd_sc_hd__dfrtp_1 c118(
.D(net64),
.RESET_B(net58),
.CLK(clk),
.Q(net65)
);

sky130_fd_sc_hd__dfrtp_2 c119(
.D(net53),
.RESET_B(net55),
.CLK(clk),
.Q(net66)
);

sky130_fd_sc_hd__and2_0 c120(
.A(net65),
.B(net63),
.X(net67)
);

sky130_fd_sc_hd__a21oi_2 c121(
.A1(net66),
.A2(net60),
.B1(net67),
.Y(net68)
);

sky130_fd_sc_hd__o31ai_1 c122(
.A1(net62),
.A2(net68),
.A3(net42),
.B1(net67),
.Y(net69)
);

sky130_fd_sc_hd__a21boi_1 c123(
.A1(net57),
.A2(net4),
.B1_N(net67),
.Y(net70)
);

sky130_fd_sc_hd__dfbbn_1 c124(
.D(net69),
.RESET_B(net11),
.SET_B(net58),
.CLK_N(clk),
.Q(out20),
.Q_N(net71)
);

sky130_fd_sc_hd__dfbbn_2 c125(
.D(net63),
.RESET_B(net69),
.SET_B(net58),
.CLK_N(clk),
.Q(out21),
.Q_N(net72)
);

sky130_fd_sc_hd__nor2b_1 c126(
.A(in20),
.B_N(in19),
.Y(net73)
);

sky130_fd_sc_hd__nand2b_1 c127(
.A_N(in19),
.B(in6),
.Y(net74)
);

sky130_fd_sc_hd__or2_4 c128(
.A(in1),
.B(in7),
.X(net75)
);

sky130_fd_sc_hd__nor2_4 c129(
.A(net73),
.B(in19),
.Y(net76)
);

sky130_fd_sc_hd__and2_1 c130(
.A(in12),
.B(in8),
.X(net77)
);

sky130_fd_sc_hd__or2b_4 c131(
.A(net77),
.B_N(in4),
.X(net78)
);

sky130_fd_sc_hd__a21o_4 c132(
.A1(in17),
.A2(in13),
.B1(net75),
.X(net79)
);

sky130_fd_sc_hd__nor2_4 c133(
.A(in4),
.B(net75),
.Y(net80)
);

sky130_fd_sc_hd__or2_4 c134(
.A(net79),
.B(in10),
.X(net81)
);

sky130_fd_sc_hd__or2b_2 c135(
.A(in8),
.B_N(net77),
.X(net82)
);

sky130_fd_sc_hd__a21oi_4 c136(
.A1(net78),
.A2(in20),
.B1(net82),
.Y(net83)
);

sky130_fd_sc_hd__nor2b_2 c137(
.A(net75),
.B_N(in0),
.Y(net84)
);

sky130_fd_sc_hd__nor2_2 c138(
.A(net82),
.B(net74),
.Y(net85)
);

sky130_fd_sc_hd__mux2_8 c139(
.A0(net80),
.A1(net82),
.S(in11),
.X(net86)
);

sky130_fd_sc_hd__and2_4 c140(
.A(in11),
.B(net84),
.X(net87)
);

sky130_fd_sc_hd__mux2_2 c141(
.A0(in0),
.A1(net85),
.S(net87),
.X(net88)
);

sky130_fd_sc_hd__or2b_1 c142(
.A(net87),
.B_N(net73),
.X(net89)
);

sky130_fd_sc_hd__or2b_4 c143(
.A(net89),
.B_N(net86),
.X(net90)
);

sky130_fd_sc_hd__o41a_1 c144(
.A1(net76),
.A2(in7),
.A3(net90),
.A4(net89),
.B1(net88),
.X(net91)
);

sky130_fd_sc_hd__or2b_4 c145(
.A(net90),
.B_N(net84),
.X(net92)
);

sky130_fd_sc_hd__nor2_2 c146(
.A(net92),
.B(net90),
.Y(net93)
);

sky130_fd_sc_hd__nor2_2 c147(
.A(in5),
.B(in38),
.Y(net94)
);

sky130_fd_sc_hd__nor2_2 c148(
.A(net94),
.B(in41),
.Y(net95)
);

sky130_fd_sc_hd__or2b_1 c149(
.A(in27),
.B_N(in13),
.X(net96)
);

sky130_fd_sc_hd__and2b_4 c150(
.A_N(in35),
.B(in13),
.X(net97)
);

sky130_fd_sc_hd__a21o_1 c151(
.A1(in37),
.A2(in5),
.B1(in23),
.X(net98)
);

sky130_fd_sc_hd__nor2_1 c152(
.A(in25),
.B(in30),
.Y(net99)
);

sky130_fd_sc_hd__nand2_4 c153(
.A(in10),
.B(in35),
.Y(net100)
);

sky130_fd_sc_hd__nor2_4 c154(
.A(in34),
.B(net100),
.Y(net101)
);

sky130_fd_sc_hd__nand2b_1 c155(
.A_N(net97),
.B(net99),
.Y(net102)
);

sky130_fd_sc_hd__or2_2 c156(
.A(net102),
.B(net101),
.X(net103)
);

sky130_fd_sc_hd__or2b_4 c157(
.A(net77),
.B_N(net73),
.X(net104)
);

sky130_fd_sc_hd__o21a_1 c158(
.A1(net96),
.A2(net81),
.B1(net102),
.X(net105)
);

sky130_fd_sc_hd__or2b_1 c159(
.A(net101),
.B_N(net102),
.X(net106)
);

sky130_fd_sc_hd__a21o_4 c160(
.A1(net84),
.A2(net96),
.B1(net75),
.X(net107)
);

sky130_fd_sc_hd__o31a_1 c161(
.A1(net106),
.A2(net100),
.A3(net97),
.B1(net102),
.X(net108)
);

sky130_fd_sc_hd__a21o_1 c162(
.A1(net100),
.A2(net108),
.B1(net102),
.X(net109)
);

sky130_fd_sc_hd__mux4_1 c163(
.A0(net108),
.A1(net102),
.A2(net109),
.A3(net103),
.S0(net104),
.S1(net106),
.X(net110)
);

sky130_fd_sc_hd__o41a_1 c164(
.A1(net97),
.A2(net106),
.A3(net110),
.A4(net109),
.B1(net94),
.X(net111)
);

sky130_fd_sc_hd__a21o_2 c165(
.A1(net105),
.A2(net108),
.B1(net101),
.X(net112)
);

sky130_fd_sc_hd__a21bo_1 c166(
.A1(net107),
.A2(net110),
.B1_N(in10),
.X(net113)
);

sky130_fd_sc_hd__and2_1 c167(
.A(net110),
.B(in35),
.X(out23)
);

sky130_fd_sc_hd__a21oi_1 c168(
.A1(in31),
.A2(net8),
.B1(in51),
.Y(net114)
);

sky130_fd_sc_hd__nor2_1 c169(
.A(net114),
.B(in9),
.Y(net115)
);

sky130_fd_sc_hd__nand2b_1 c170(
.A_N(in32),
.B(net83),
.Y(net116)
);

sky130_fd_sc_hd__o21a_1 c171(
.A1(net2),
.A2(net115),
.B1(net10),
.X(net117)
);

sky130_fd_sc_hd__o21bai_1 c172(
.A1(net80),
.A2(net114),
.B1_N(in51),
.Y(net118)
);

sky130_fd_sc_hd__and2b_1 c173(
.A_N(net8),
.B(out23),
.X(net119)
);

sky130_fd_sc_hd__nor2b_1 c174(
.A(net116),
.B_N(in51),
.Y(net120)
);

sky130_fd_sc_hd__nand2_4 c175(
.A(net10),
.B(in7),
.Y(net121)
);

sky130_fd_sc_hd__and2_2 c176(
.A(net121),
.B(net119),
.X(out30)
);

sky130_fd_sc_hd__or2_2 c177(
.A(net115),
.B(in51),
.X(net122)
);

sky130_fd_sc_hd__and2b_2 c178(
.A_N(net89),
.B(net114),
.X(net123)
);

sky130_fd_sc_hd__nand2_1 c179(
.A(net123),
.B(net103),
.Y(net124)
);

sky130_fd_sc_hd__mux2_1 c180(
.A0(in29),
.A1(net124),
.S(in51),
.X(net125)
);

sky130_fd_sc_hd__o21a_1 c181(
.A1(net121),
.A2(net83),
.B1(net119),
.X(net126)
);

sky130_fd_sc_hd__nor2_2 c182(
.A(net120),
.B(in51),
.Y(net127)
);

sky130_fd_sc_hd__and2_2 c183(
.A(net92),
.B(in51),
.X(net128)
);

sky130_fd_sc_hd__nor2b_4 c184(
.A(net128),
.B_N(net123),
.Y(net129)
);

sky130_fd_sc_hd__a21o_2 c185(
.A1(in48),
.A2(net121),
.B1(net129),
.X(net130)
);

sky130_fd_sc_hd__nor2b_2 c186(
.A(net125),
.B_N(net129),
.Y(net131)
);

sky130_fd_sc_hd__o21bai_4 c187(
.A1(net129),
.A2(net131),
.B1_N(net130),
.Y(net132)
);

sky130_fd_sc_hd__o31ai_4 c188(
.A1(net122),
.A2(net132),
.A3(net128),
.B1(net119),
.Y(net133)
);

sky130_fd_sc_hd__or2b_4 c189(
.A(in30),
.B_N(net116),
.X(net134)
);

sky130_fd_sc_hd__and2b_2 c190(
.A_N(net101),
.B(in30),
.X(net135)
);

sky130_fd_sc_hd__and2b_4 c191(
.A_N(net130),
.B(in38),
.X(net136)
);

sky130_fd_sc_hd__nand2_2 c192(
.A(net134),
.B(net135),
.Y(net137)
);

sky130_fd_sc_hd__or2_2 c193(
.A(net120),
.B(net29),
.X(out41)
);

sky130_fd_sc_hd__a21o_2 c194(
.A1(net136),
.A2(net134),
.B1(net83),
.X(net138)
);

sky130_fd_sc_hd__a21boi_1 c195(
.A1(net23),
.A2(net119),
.B1_N(net27),
.Y(net139)
);

sky130_fd_sc_hd__o41a_2 c196(
.A1(net12),
.A2(net137),
.A3(net134),
.A4(net118),
.B1(net99),
.X(net140)
);

sky130_fd_sc_hd__and2b_1 c197(
.A_N(in50),
.B(in13),
.X(net141)
);

sky130_fd_sc_hd__nand2b_2 c198(
.A_N(net27),
.B(net139),
.Y(net142)
);

sky130_fd_sc_hd__nor2b_4 c199(
.A(net83),
.B_N(net140),
.Y(net143)
);

sky130_fd_sc_hd__o41a_4 c200(
.A1(net137),
.A2(net139),
.A3(net143),
.A4(net141),
.B1(net142),
.X(net144)
);

sky130_fd_sc_hd__nand2b_2 c201(
.A_N(net133),
.B(net142),
.Y(net145)
);

sky130_fd_sc_hd__and2_1 c202(
.A(net145),
.B(net141),
.X(net146)
);

sky130_fd_sc_hd__and2_4 c203(
.A(net143),
.B(net138),
.X(net147)
);

sky130_fd_sc_hd__or2b_4 c204(
.A(net139),
.B_N(net142),
.X(net148)
);

sky130_fd_sc_hd__nor2_4 c205(
.A(net17),
.B(net137),
.Y(net149)
);

sky130_fd_sc_hd__mux2_8 c206(
.A0(net149),
.A1(net141),
.S(net112),
.X(net150)
);

sky130_fd_sc_hd__mux4_4 c207(
.A0(net146),
.A1(net136),
.A2(net149),
.A3(net150),
.S0(net114),
.S1(net138),
.X(net151)
);

sky130_fd_sc_hd__mux4_1 c208(
.A0(net134),
.A1(net140),
.A2(in15),
.A3(net149),
.S0(net142),
.S1(net151),
.X(net152)
);

sky130_fd_sc_hd__a21oi_2 c209(
.A1(net151),
.A2(net150),
.B1(net147),
.Y(net153)
);

sky130_fd_sc_hd__nand2_2 c210(
.A(net49),
.B(net148),
.Y(net154)
);

sky130_fd_sc_hd__nor2b_1 c211(
.A(net33),
.B_N(net50),
.Y(net155)
);

sky130_fd_sc_hd__nor2b_2 c212(
.A(net147),
.B_N(net150),
.Y(out40)
);

sky130_fd_sc_hd__and2_0 c213(
.A(net116),
.B(net144),
.X(net156)
);

sky130_fd_sc_hd__a21o_1 c214(
.A1(net39),
.A2(net12),
.B1(net147),
.X(net157)
);

sky130_fd_sc_hd__inv_8 c215(
.A(net639),
.Y(net158)
);

sky130_fd_sc_hd__and2b_2 c216(
.A_N(net50),
.B(in51),
.X(net159)
);

sky130_fd_sc_hd__clkinv_4 c217(
.A(net638),
.Y(net160)
);

sky130_fd_sc_hd__and2b_1 c218(
.A_N(net158),
.B(net160),
.X(out31)
);

sky130_fd_sc_hd__nand2b_1 c219(
.A_N(net160),
.B(net158),
.Y(net161)
);

sky130_fd_sc_hd__sdfrbp_1 c220(
.D(net40),
.RESET_B(net152),
.SCD(net160),
.SCE(out31),
.CLK(clk),
.Q(net163),
.Q_N(net162)
);

sky130_fd_sc_hd__a21bo_1 c221(
.A1(net15),
.A2(net142),
.B1_N(net157),
.X(out28)
);

sky130_fd_sc_hd__nand2b_1 c222(
.A_N(net161),
.B(out28),
.Y(net164)
);

sky130_fd_sc_hd__mux4_1 c223(
.A0(net150),
.A1(net141),
.A2(net160),
.A3(net114),
.S0(out28),
.S1(net157),
.X(net165)
);

sky130_fd_sc_hd__or2b_4 c224(
.A(net142),
.B_N(net155),
.X(net166)
);

sky130_fd_sc_hd__dfbbp_1 c225(
.D(net119),
.RESET_B(net162),
.SET_B(net165),
.CLK(clk),
.Q(net168),
.Q_N(net167)
);

sky130_fd_sc_hd__sdfxbp_1 c226(
.D(net165),
.SCD(net167),
.SCE(out31),
.CLK(clk),
.Q(net170),
.Q_N(net169)
);

sky130_fd_sc_hd__mux4_1 c227(
.A0(net43),
.A1(out31),
.A2(net116),
.A3(net42),
.S0(out30),
.S1(net159),
.X(net171)
);

sky130_fd_sc_hd__nand2_4 c228(
.A(net168),
.B(net39),
.Y(net172)
);

sky130_fd_sc_hd__mux4_4 c229(
.A0(net171),
.A1(net172),
.A2(net47),
.A3(net164),
.S0(net33),
.S1(out31),
.X(net173)
);

sky130_fd_sc_hd__mux4_4 c230(
.A0(net159),
.A1(net169),
.A2(net172),
.A3(out31),
.S0(in14),
.S1(net644),
.X(net174)
);

sky130_fd_sc_hd__o21bai_2 c231(
.A1(net148),
.A2(net46),
.B1_N(net79),
.Y(net175)
);

sky130_fd_sc_hd__and2_4 c232(
.A(net86),
.B(net46),
.X(net176)
);

sky130_fd_sc_hd__dfrtp_4 c233(
.D(net174),
.RESET_B(net67),
.CLK(clk),
.Q(net177)
);

sky130_fd_sc_hd__mux2_1 c234(
.A0(net176),
.A1(net67),
.S(net47),
.X(out9)
);

sky130_fd_sc_hd__sdfxbp_2 c235(
.D(net52),
.SCD(in51),
.SCE(out9),
.CLK(clk),
.Q(net179),
.Q_N(net178)
);

sky130_fd_sc_hd__dfsbp_1 c236(
.D(net140),
.SET_B(net174),
.CLK(clk),
.Q(net181),
.Q_N(net180)
);

sky130_fd_sc_hd__or2_4 c237(
.A(net82),
.B(net112),
.X(net182)
);

sky130_fd_sc_hd__nor2b_1 c238(
.A(net181),
.B_N(net175),
.Y(net183)
);

sky130_fd_sc_hd__nand2b_2 c239(
.A_N(net182),
.B(net176),
.Y(net184)
);

sky130_fd_sc_hd__and2b_1 c240(
.A_N(net177),
.B(out21),
.X(net185)
);

sky130_fd_sc_hd__nor2_1 c241(
.A(net185),
.B(net47),
.Y(out0)
);

sky130_fd_sc_hd__or2_1 c242(
.A(net42),
.B(out40),
.X(net186)
);

sky130_fd_sc_hd__mux4_1 c243(
.A0(net59),
.A1(net154),
.A2(out0),
.A3(net46),
.S0(net178),
.S1(out9),
.X(net187)
);

sky130_fd_sc_hd__o21ai_2 c244(
.A1(net185),
.A2(net182),
.B1(net646),
.Y(net188)
);

sky130_fd_sc_hd__sdfxtp_1 c245(
.D(net70),
.SCD(net180),
.SCE(out9),
.CLK(clk),
.Q(net189)
);

sky130_fd_sc_hd__sdfxtp_2 c246(
.D(net179),
.SCD(net186),
.SCE(net183),
.CLK(clk),
.Q(out24)
);

sky130_fd_sc_hd__sdfrbp_2 c247(
.D(net188),
.RESET_B(net184),
.SCD(net189),
.SCE(out24),
.CLK(clk),
.Q(net191),
.Q_N(net190)
);

sky130_fd_sc_hd__o21bai_1 c248(
.A1(net175),
.A2(net185),
.B1_N(net70),
.Y(net192)
);

sky130_fd_sc_hd__mux4_1 c249(
.A0(net189),
.A1(out6),
.A2(net190),
.A3(out30),
.S0(out31),
.S1(out9),
.X(net193)
);

sky130_fd_sc_hd__sdfxtp_4 c250(
.D(out9),
.SCD(net148),
.SCE(net647),
.CLK(clk),
.Q(net194)
);

sky130_fd_sc_hd__a21boi_2 c251(
.A1(net191),
.A2(net194),
.B1_N(net647),
.Y(out22)
);

sky130_fd_sc_hd__nand2b_2 c252(
.A_N(net91),
.B(in6),
.Y(net195)
);

sky130_fd_sc_hd__clkbuf_4 c253(
.A(net73),
.X(net196)
);

sky130_fd_sc_hd__and2b_2 c254(
.A_N(in14),
.B(net87),
.X(net197)
);

sky130_fd_sc_hd__and2_2 c255(
.A(net197),
.B(net91),
.X(net198)
);

sky130_fd_sc_hd__inv_1 c256(
.A(net78),
.Y(net199)
);

sky130_fd_sc_hd__clkinv_2 c257(
.A(in12),
.Y(net200)
);

sky130_fd_sc_hd__or2_2 c258(
.A(net200),
.B(net88),
.X(net201)
);

sky130_fd_sc_hd__or2_1 c259(
.A(net201),
.B(net200),
.X(net202)
);

sky130_fd_sc_hd__nor2b_2 c260(
.A(net198),
.B_N(net201),
.Y(net203)
);

sky130_fd_sc_hd__nand2_1 c261(
.A(net202),
.B(net200),
.Y(net204)
);

sky130_fd_sc_hd__or2_2 c262(
.A(net203),
.B(net201),
.X(net205)
);

sky130_fd_sc_hd__nor2b_1 c263(
.A(net85),
.B_N(net78),
.Y(net206)
);

sky130_fd_sc_hd__and2_1 c264(
.A(net205),
.B(net206),
.X(net207)
);

sky130_fd_sc_hd__or2_1 c265(
.A(net204),
.B(net202),
.X(net208)
);

sky130_fd_sc_hd__nor2_1 c266(
.A(net199),
.B(net208),
.Y(net209)
);

sky130_fd_sc_hd__and2_4 c267(
.A(net202),
.B(net204),
.X(net210)
);

sky130_fd_sc_hd__nand2b_2 c268(
.A_N(net195),
.B(net196),
.Y(net211)
);

sky130_fd_sc_hd__nand2_4 c269(
.A(net206),
.B(net210),
.Y(net212)
);

sky130_fd_sc_hd__o21ai_4 c270(
.A1(net210),
.A2(net200),
.B1(net211),
.Y(net213)
);

sky130_fd_sc_hd__or2_1 c271(
.A(net212),
.B(net213),
.X(net214)
);

sky130_fd_sc_hd__o21bai_1 c272(
.A1(net213),
.A2(net211),
.B1_N(net214),
.Y(net215)
);

sky130_fd_sc_hd__or2_2 c273(
.A(in28),
.B(in40),
.X(net216)
);

sky130_fd_sc_hd__a21boi_4 c274(
.A1(net203),
.A2(net81),
.B1_N(net216),
.Y(net217)
);

sky130_fd_sc_hd__or2_2 c275(
.A(in26),
.B(net95),
.X(net218)
);

sky130_fd_sc_hd__nor2b_4 c276(
.A(net207),
.B_N(net216),
.Y(net219)
);

sky130_fd_sc_hd__and2_1 c277(
.A(in1),
.B(net200),
.X(net220)
);

sky130_fd_sc_hd__or2b_4 c278(
.A(in33),
.B_N(net98),
.X(net221)
);

sky130_fd_sc_hd__nor2_2 c279(
.A(net221),
.B(net220),
.Y(net222)
);

sky130_fd_sc_hd__and2b_4 c280(
.A_N(net214),
.B(net113),
.X(net223)
);

sky130_fd_sc_hd__or2b_2 c281(
.A(net220),
.B_N(net88),
.X(net224)
);

sky130_fd_sc_hd__and2_4 c282(
.A(net219),
.B(net223),
.X(net225)
);

sky130_fd_sc_hd__nor2b_1 c283(
.A(net222),
.B_N(net109),
.Y(net226)
);

sky130_fd_sc_hd__nor2_2 c284(
.A(net81),
.B(net222),
.Y(net227)
);

sky130_fd_sc_hd__or2_2 c285(
.A(net217),
.B(net81),
.X(net228)
);

sky130_fd_sc_hd__o31a_2 c286(
.A1(net219),
.A2(net207),
.A3(net227),
.B1(net224),
.X(net229)
);

sky130_fd_sc_hd__nand2_2 c287(
.A(net229),
.B(net224),
.Y(net230)
);

sky130_fd_sc_hd__o31ai_2 c288(
.A1(net227),
.A2(net214),
.A3(net230),
.B1(net224),
.Y(net231)
);

sky130_fd_sc_hd__and2_4 c289(
.A(net227),
.B(net225),
.X(net232)
);

sky130_fd_sc_hd__o21bai_1 c290(
.A1(net231),
.A2(net230),
.B1_N(net225),
.Y(net233)
);

sky130_fd_sc_hd__sdfbbn_1 c291(
.D(net226),
.RESET_B(out23),
.SCD(net233),
.SCE(net225),
.SET_B(net98),
.CLK_N(clk),
.Q(net235),
.Q_N(net234)
);

sky130_fd_sc_hd__and2_4 c292(
.A(net197),
.B(net224),
.X(net236)
);

sky130_fd_sc_hd__dfsbp_2 c293(
.D(net233),
.SET_B(net236),
.CLK(clk),
.Q(net238),
.Q_N(net237)
);

sky130_fd_sc_hd__nor2_4 c294(
.A(in9),
.B(net225),
.Y(net239)
);

sky130_fd_sc_hd__o21ba_2 c295(
.A1(net126),
.A2(net223),
.B1_N(net88),
.X(net240)
);

sky130_fd_sc_hd__and2b_4 c296(
.A_N(net239),
.B(net131),
.X(net241)
);

sky130_fd_sc_hd__nand2b_4 c297(
.A_N(net240),
.B(net225),
.Y(net242)
);

sky130_fd_sc_hd__nor2_1 c298(
.A(net128),
.B(net126),
.Y(net243)
);

sky130_fd_sc_hd__or2b_1 c299(
.A(net200),
.B_N(net242),
.X(net244)
);

sky130_fd_sc_hd__nor2_2 c300(
.A(net241),
.B(net118),
.Y(net245)
);

sky130_fd_sc_hd__and2_0 c301(
.A(net222),
.B(net200),
.X(net246)
);

sky130_fd_sc_hd__or2_4 c302(
.A(net131),
.B(net242),
.X(net247)
);

sky130_fd_sc_hd__nand2_1 c303(
.A(net123),
.B(net223),
.Y(net248)
);

sky130_fd_sc_hd__and2_0 c304(
.A(net230),
.B(net242),
.X(net249)
);

sky130_fd_sc_hd__and2_0 c305(
.A(net223),
.B(net200),
.X(net250)
);

sky130_fd_sc_hd__a21oi_1 c306(
.A1(net246),
.A2(net249),
.B1(net126),
.Y(net251)
);

sky130_fd_sc_hd__and2_1 c307(
.A(net247),
.B(net100),
.X(net252)
);

sky130_fd_sc_hd__nand2_2 c308(
.A(net250),
.B(net240),
.Y(out45)
);

sky130_fd_sc_hd__mux4_4 c309(
.A0(net243),
.A1(net200),
.A2(net252),
.A3(net245),
.S0(in23),
.S1(net223),
.X(net253)
);

sky130_fd_sc_hd__nand2_1 c310(
.A(net244),
.B(net247),
.Y(net254)
);

sky130_fd_sc_hd__nand2_2 c311(
.A(net129),
.B(out45),
.Y(net255)
);

sky130_fd_sc_hd__dfstp_1 c312(
.D(net251),
.SET_B(net222),
.CLK(clk),
.Q(net256)
);

sky130_fd_sc_hd__mux4_2 c313(
.A0(net256),
.A1(net249),
.A2(net251),
.A3(net240),
.S0(net252),
.S1(net648),
.X(net257)
);

sky130_fd_sc_hd__dfstp_2 c314(
.D(net251),
.SET_B(net649),
.CLK(clk),
.Q(net258)
);

sky130_fd_sc_hd__nand2b_1 c315(
.A_N(net248),
.B(net138),
.Y(net259)
);

sky130_fd_sc_hd__o31a_2 c316(
.A1(in43),
.A2(net114),
.A3(net258),
.B1(in51),
.X(net260)
);

sky130_fd_sc_hd__nor2_4 c317(
.A(net220),
.B(net648),
.Y(out29)
);

sky130_fd_sc_hd__mux2_8 c318(
.A0(in40),
.A1(net114),
.S(in23),
.X(net261)
);

sky130_fd_sc_hd__nand2b_2 c319(
.A_N(net260),
.B(out29),
.Y(net262)
);

sky130_fd_sc_hd__dfbbn_1 c320(
.D(net153),
.RESET_B(net95),
.SET_B(net225),
.CLK_N(clk),
.Q(net264),
.Q_N(net263)
);

sky130_fd_sc_hd__o21ai_4 c321(
.A1(net138),
.A2(net225),
.B1(net263),
.Y(net265)
);

sky130_fd_sc_hd__a21bo_2 c322(
.A1(in19),
.A2(net263),
.B1_N(net258),
.X(net266)
);

sky130_fd_sc_hd__o21ai_4 c323(
.A1(net266),
.A2(net24),
.B1(net247),
.Y(net267)
);

sky130_fd_sc_hd__mux4_1 c324(
.A0(net74),
.A1(net267),
.A2(net259),
.A3(net138),
.S0(in38),
.S1(net648),
.X(net268)
);

sky130_fd_sc_hd__mux4_4 c325(
.A0(net1),
.A1(net264),
.A2(out45),
.A3(net204),
.S0(out29),
.S1(net650),
.X(net269)
);

sky130_fd_sc_hd__and2b_2 c326(
.A_N(net269),
.B(out11),
.X(net270)
);

sky130_fd_sc_hd__and2_4 c327(
.A(net261),
.B(out29),
.X(net271)
);

sky130_fd_sc_hd__nand2_4 c328(
.A(net271),
.B(net259),
.Y(out51)
);

sky130_fd_sc_hd__dfbbn_2 c329(
.D(net270),
.RESET_B(net247),
.SET_B(out51),
.CLK_N(clk),
.Q(net272)
);

sky130_fd_sc_hd__o21ba_2 c330(
.A1(net264),
.A2(net269),
.B1_N(net265),
.X(net273)
);

sky130_fd_sc_hd__o21ba_1 c331(
.A1(net262),
.A2(net264),
.B1_N(out51),
.X(net274)
);

sky130_fd_sc_hd__dfbbp_1 c332(
.D(in7),
.RESET_B(net270),
.SET_B(net267),
.CLK(clk),
.Q(net276),
.Q_N(net275)
);

sky130_fd_sc_hd__dfstp_4 c333(
.D(net274),
.SET_B(net650),
.CLK(clk),
.Q(out8)
);

sky130_fd_sc_hd__a21bo_1 c334(
.A1(net272),
.A2(out8),
.B1_N(out51),
.X(net277)
);

sky130_fd_sc_hd__mux4_2 c335(
.A0(net274),
.A1(net21),
.A2(net204),
.A3(out51),
.S0(net144),
.S1(net270),
.X(net278)
);

sky130_fd_sc_hd__dlrbn_1 c336(
.D(net164),
.RESET_B(net112),
.GATE_N(clk),
.Q(net280),
.Q_N(net279)
);

sky130_fd_sc_hd__nand2b_4 c337(
.A_N(net163),
.B(net204),
.Y(net281)
);

sky130_fd_sc_hd__and2b_2 c338(
.A_N(net172),
.B(net279),
.X(net282)
);

sky130_fd_sc_hd__and2_1 c339(
.A(net170),
.B(net104),
.X(net283)
);

sky130_fd_sc_hd__or2b_4 c340(
.A(net31),
.B_N(net144),
.X(net284)
);

sky130_fd_sc_hd__and2_0 c341(
.A(net144),
.B(net118),
.X(net285)
);

sky130_fd_sc_hd__sdfxbp_1 c342(
.D(net284),
.SCD(net265),
.SCE(net164),
.CLK(clk),
.Q(net286)
);

sky130_fd_sc_hd__nand2_1 c343(
.A(net285),
.B(net74),
.Y(net287)
);

sky130_fd_sc_hd__nor2b_4 c344(
.A(net225),
.B_N(out28),
.Y(net288)
);

sky130_fd_sc_hd__nor2_4 c345(
.A(net156),
.B(net287),
.Y(net289)
);

sky130_fd_sc_hd__and2b_4 c346(
.A_N(net289),
.B(net281),
.X(net290)
);

sky130_fd_sc_hd__and2b_4 c347(
.A_N(net157),
.B(net209),
.X(net291)
);

sky130_fd_sc_hd__and2_0 c348(
.A(net45),
.B(net225),
.X(net292)
);

sky130_fd_sc_hd__o31ai_1 c349(
.A1(net280),
.A2(net48),
.A3(net38),
.B1(net225),
.Y(net293)
);

sky130_fd_sc_hd__sdfbbn_2 c350(
.D(net293),
.RESET_B(net288),
.SCD(net156),
.SCE(out8),
.SET_B(out29),
.CLK_N(clk),
.Q(net294)
);

sky130_fd_sc_hd__dlrbn_2 c351(
.D(net288),
.RESET_B(net45),
.GATE_N(clk),
.Q(net296),
.Q_N(net295)
);

sky130_fd_sc_hd__nor2b_2 c352(
.A(net294),
.B_N(net296),
.Y(net297)
);

sky130_fd_sc_hd__o41a_1 c353(
.A1(net291),
.A2(net161),
.A3(out11),
.A4(net295),
.B1(net46),
.X(net298)
);

sky130_fd_sc_hd__sdfxbp_2 c354(
.D(net282),
.SCD(net298),
.SCE(net161),
.CLK(clk),
.Q(net300),
.Q_N(net299)
);

sky130_fd_sc_hd__sdfxtp_1 c355(
.D(net286),
.SCD(net297),
.SCE(net298),
.CLK(clk),
.Q(net301)
);

sky130_fd_sc_hd__mux4_4 c356(
.A0(net301),
.A1(net225),
.A2(net295),
.A3(net291),
.S0(net284),
.S1(out8),
.X(net302)
);

sky130_fd_sc_hd__a21boi_0 c357(
.A1(net283),
.A2(net104),
.B1_N(out45),
.Y(net303)
);

sky130_fd_sc_hd__a21boi_2 c358(
.A1(net259),
.A2(net296),
.B1_N(out24),
.Y(net304)
);

sky130_fd_sc_hd__sdfxtp_2 c359(
.D(net48),
.SCD(net298),
.SCE(net60),
.CLK(clk),
.Q(net305)
);

sky130_fd_sc_hd__dlrbp_1 c360(
.D(net183),
.RESET_B(out31),
.GATE(clk),
.Q(net307),
.Q_N(net306)
);

sky130_fd_sc_hd__dlrbp_2 c361(
.D(net184),
.RESET_B(net177),
.GATE(clk),
.Q(net308)
);

sky130_fd_sc_hd__dlrtn_1 c362(
.D(net192),
.RESET_B(net305),
.GATE_N(clk),
.Q(net309)
);

sky130_fd_sc_hd__a21oi_2 c363(
.A1(net68),
.A2(net303),
.B1(net295),
.Y(net310)
);

sky130_fd_sc_hd__nor2_4 c364(
.A(net305),
.B(net71),
.Y(net311)
);

sky130_fd_sc_hd__a21bo_1 c365(
.A1(net308),
.A2(net61),
.B1_N(net306),
.X(net312)
);

sky130_fd_sc_hd__sdfxtp_4 c366(
.D(net154),
.SCD(out9),
.SCE(in51),
.CLK(clk),
.Q(out44)
);

sky130_fd_sc_hd__a21boi_1 c367(
.A1(in13),
.A2(net194),
.B1_N(in51),
.Y(net313)
);

sky130_fd_sc_hd__a21boi_1 c368(
.A1(in51),
.A2(net311),
.B1_N(out41),
.Y(net314)
);

sky130_fd_sc_hd__dfbbn_1 c369(
.D(net67),
.RESET_B(net310),
.SET_B(net61),
.CLK_N(clk),
.Q(net315)
);

sky130_fd_sc_hd__o21bai_2 c370(
.A1(net61),
.A2(net305),
.B1_N(out24),
.Y(net316)
);

sky130_fd_sc_hd__dlrtn_2 c371(
.D(net58),
.RESET_B(net316),
.GATE_N(clk),
.Q(net317)
);

sky130_fd_sc_hd__or2b_4 c372(
.A(net292),
.B_N(net315),
.X(out43)
);

sky130_fd_sc_hd__o21bai_4 c373(
.A1(net112),
.A2(net317),
.B1_N(out45),
.Y(net318)
);

sky130_fd_sc_hd__o31a_2 c374(
.A1(net314),
.A2(net318),
.A3(out21),
.B1(net209),
.X(net319)
);

sky130_fd_sc_hd__sdfrtn_1 c375(
.D(net319),
.RESET_B(net312),
.SCD(out31),
.SCE(out44),
.CLK_N(clk),
.Q(net320)
);

sky130_fd_sc_hd__dfbbn_2 c376(
.D(net313),
.RESET_B(net320),
.SET_B(net319),
.CLK_N(clk),
.Q(net322),
.Q_N(net321)
);

sky130_fd_sc_hd__o31ai_2 c377(
.A1(net317),
.A2(net318),
.A3(out0),
.B1(net316),
.Y(out35)
);

sky130_fd_sc_hd__or2_2 c378(
.A(net215),
.B(net198),
.X(net323)
);

sky130_fd_sc_hd__and2_2 c379(
.A(in17),
.B(net211),
.X(net324)
);

sky130_fd_sc_hd__nor2_1 c380(
.A(net211),
.B(net215),
.Y(net325)
);

sky130_fd_sc_hd__nand2b_2 c381(
.A_N(net90),
.B(net93),
.Y(net326)
);

sky130_fd_sc_hd__and2_0 c382(
.A(net326),
.B(net79),
.X(net327)
);

sky130_fd_sc_hd__and2_0 c383(
.A(net323),
.B(net326),
.X(net328)
);

sky130_fd_sc_hd__and2_1 c384(
.A(net327),
.B(net326),
.X(net329)
);

sky130_fd_sc_hd__and2_4 c385(
.A(net323),
.B(in15),
.X(net330)
);

sky130_fd_sc_hd__or2b_2 c386(
.A(net329),
.B_N(net330),
.X(net331)
);

sky130_fd_sc_hd__or2_2 c387(
.A(net330),
.B(net328),
.X(net332)
);

sky130_fd_sc_hd__clkinv_1 c388(
.A(net196),
.Y(net333)
);

sky130_fd_sc_hd__nor2b_4 c389(
.A(net333),
.B_N(net332),
.Y(net334)
);

sky130_fd_sc_hd__mux2_4 c390(
.A0(net327),
.A1(net324),
.S(net211),
.X(net335)
);

sky130_fd_sc_hd__and2_4 c391(
.A(net331),
.B(net196),
.X(net336)
);

sky130_fd_sc_hd__and2b_4 c392(
.A_N(net325),
.B(net333),
.X(net337)
);

sky130_fd_sc_hd__and2_2 c393(
.A(net331),
.B(net332),
.X(net338)
);

sky130_fd_sc_hd__nor2_1 c394(
.A(net335),
.B(net328),
.Y(net339)
);

sky130_fd_sc_hd__sdfbbp_1 c395(
.D(net330),
.RESET_B(net336),
.SCD(net338),
.SCE(net339),
.SET_B(net333),
.CLK(clk),
.Q(net341),
.Q_N(net340)
);

sky130_fd_sc_hd__dlrtn_4 c396(
.D(net334),
.RESET_B(net340),
.GATE_N(clk),
.Q(net342)
);

sky130_fd_sc_hd__dlrtp_1 c397(
.D(net338),
.RESET_B(net330),
.GATE(clk),
.Q(net343)
);

sky130_fd_sc_hd__or2_1 c398(
.A(net341),
.B(net328),
.X(out39)
);

sky130_fd_sc_hd__and2b_4 c399(
.A_N(net235),
.B(net104),
.X(net344)
);

sky130_fd_sc_hd__and2_2 c400(
.A(net208),
.B(out39),
.X(net345)
);

sky130_fd_sc_hd__nand2_4 c401(
.A(net236),
.B(net237),
.Y(net346)
);

sky130_fd_sc_hd__and2b_2 c402(
.A_N(net342),
.B(net226),
.X(net347)
);

sky130_fd_sc_hd__or2_1 c403(
.A(net218),
.B(net346),
.X(out4)
);

sky130_fd_sc_hd__dlrtp_2 c404(
.D(net344),
.RESET_B(net345),
.GATE(clk),
.Q(net348)
);

sky130_fd_sc_hd__dlrtp_4 c405(
.D(net224),
.RESET_B(net345),
.GATE(clk),
.Q(net349)
);

sky130_fd_sc_hd__dfbbp_1 c406(
.D(net345),
.RESET_B(net234),
.SET_B(net343),
.CLK(clk),
.Q(net351),
.Q_N(net350)
);

sky130_fd_sc_hd__and2b_1 c407(
.A_N(net348),
.B(net195),
.X(net352)
);

sky130_fd_sc_hd__or2_1 c408(
.A(net109),
.B(out4),
.X(net353)
);

sky130_fd_sc_hd__a21bo_2 c409(
.A1(net75),
.A2(net353),
.B1_N(net347),
.X(net354)
);

sky130_fd_sc_hd__and2_4 c410(
.A(net98),
.B(net350),
.X(net355)
);

sky130_fd_sc_hd__and2_1 c411(
.A(net353),
.B(net347),
.X(net356)
);

sky130_fd_sc_hd__nand2b_2 c412(
.A_N(net346),
.B(net344),
.Y(net357)
);

sky130_fd_sc_hd__mux2_8 c413(
.A0(net351),
.A1(net226),
.S(net216),
.X(net358)
);

sky130_fd_sc_hd__o41a_1 c414(
.A1(net358),
.A2(net351),
.A3(net352),
.A4(net353),
.B1(out4),
.X(net359)
);

sky130_fd_sc_hd__edfxbp_1 c415(
.D(net336),
.DE(net356),
.CLK(clk),
.Q(net361),
.Q_N(net360)
);

sky130_fd_sc_hd__nor2_2 c416(
.A(net228),
.B(net359),
.Y(net362)
);

sky130_fd_sc_hd__o21bai_4 c417(
.A1(net356),
.A2(net353),
.B1_N(net357),
.Y(net363)
);

sky130_fd_sc_hd__sdfbbn_1 c418(
.D(net349),
.RESET_B(net345),
.SCD(net342),
.SCE(net358),
.SET_B(out4),
.CLK_N(clk),
.Q(net364)
);

sky130_fd_sc_hd__o21ba_2 c419(
.A1(net357),
.A2(net364),
.B1_N(net358),
.X(net365)
);

sky130_fd_sc_hd__a21boi_2 c420(
.A1(net353),
.A2(net359),
.B1_N(net242),
.Y(net366)
);

sky130_fd_sc_hd__a21o_2 c421(
.A1(in38),
.A2(net220),
.B1(net359),
.X(net367)
);

sky130_fd_sc_hd__a21bo_1 c422(
.A1(net357),
.A2(net355),
.B1_N(in38),
.X(net368)
);

sky130_fd_sc_hd__or2_4 c423(
.A(in18),
.B(net220),
.X(net369)
);

sky130_fd_sc_hd__edfxtp_1 c424(
.D(net254),
.DE(net220),
.CLK(clk),
.Q(net370)
);

sky130_fd_sc_hd__sdlclkp_1 c425(
.GATE(net245),
.SCE(net103),
.CLK(clk),
.GCLK(net371)
);

sky130_fd_sc_hd__nand2_2 c426(
.A(net240),
.B(net99),
.Y(net372)
);

sky130_fd_sc_hd__or2b_1 c427(
.A(net362),
.B_N(net371),
.X(net373)
);

sky130_fd_sc_hd__a21oi_2 c428(
.A1(net373),
.A2(net371),
.B1(net367),
.Y(net374)
);

sky130_fd_sc_hd__or2_1 c429(
.A(net249),
.B(net368),
.X(net375)
);

sky130_fd_sc_hd__o21ba_4 c430(
.A1(net365),
.A2(net117),
.B1_N(net362),
.X(net376)
);

sky130_fd_sc_hd__or2_4 c431(
.A(net374),
.B(net361),
.X(net377)
);

sky130_fd_sc_hd__and2b_4 c432(
.A_N(net366),
.B(net359),
.X(net378)
);

sky130_fd_sc_hd__sdfxbp_1 c433(
.D(net374),
.SCD(net348),
.SCE(net378),
.CLK(clk),
.Q(net380),
.Q_N(net379)
);

sky130_fd_sc_hd__o21ba_4 c434(
.A1(net370),
.A2(net195),
.B1_N(net369),
.X(out32)
);

sky130_fd_sc_hd__o21ai_2 c435(
.A1(net373),
.A2(net356),
.B1(net370),
.Y(net381)
);

sky130_fd_sc_hd__sdfbbn_2 c436(
.D(net88),
.RESET_B(net378),
.SCD(net375),
.SCE(net353),
.SET_B(net381),
.CLK_N(clk),
.Q(net383),
.Q_N(net382)
);

sky130_fd_sc_hd__o41a_2 c437(
.A1(net368),
.A2(in41),
.A3(net383),
.A4(net374),
.B1(net367),
.X(net384)
);

sky130_fd_sc_hd__a21boi_2 c438(
.A1(net380),
.A2(net384),
.B1_N(net383),
.Y(net385)
);

sky130_fd_sc_hd__sdfrtp_1 c439(
.D(net385),
.RESET_B(net371),
.SCD(net379),
.SCE(net384),
.CLK(clk),
.Q(net386)
);

sky130_fd_sc_hd__sdfxbp_2 c440(
.D(net255),
.SCD(net385),
.SCE(net381),
.CLK(clk),
.Q(net387)
);

sky130_fd_sc_hd__sdlclkp_2 c441(
.GATE(net258),
.SCE(net277),
.CLK(clk),
.GCLK(net388)
);

sky130_fd_sc_hd__sdlclkp_4 c442(
.GATE(net265),
.SCE(net375),
.CLK(clk),
.GCLK(net389)
);

sky130_fd_sc_hd__nand2_1 c443(
.A(in15),
.B(net381),
.Y(net390)
);

sky130_fd_sc_hd__or2b_2 c444(
.A(net29),
.B_N(out8),
.X(net391)
);

sky130_fd_sc_hd__nand2b_4 c445(
.A_N(net386),
.B(net24),
.Y(net392)
);

sky130_fd_sc_hd__nand2b_4 c446(
.A_N(net387),
.B(net391),
.Y(net393)
);

sky130_fd_sc_hd__nand2_2 c447(
.A(net393),
.B(net363),
.Y(net394)
);

sky130_fd_sc_hd__sdfbbp_1 c448(
.D(net394),
.RESET_B(out41),
.SCD(net220),
.SCE(net252),
.SET_B(net391),
.CLK(clk),
.Q(net396),
.Q_N(net395)
);

sky130_fd_sc_hd__o21ai_0 c449(
.A1(net276),
.A2(net339),
.B1(net145),
.Y(net397)
);

sky130_fd_sc_hd__nor2_2 c450(
.A(net391),
.B(net651),
.Y(net398)
);

sky130_fd_sc_hd__sdfrtp_2 c451(
.D(net397),
.RESET_B(net274),
.SCD(net275),
.SCE(net391),
.CLK(clk),
.Q(out19)
);

sky130_fd_sc_hd__sdfrtp_4 c452(
.D(net376),
.RESET_B(net252),
.SCD(net394),
.SCE(net28),
.CLK(clk),
.Q(net399)
);

sky130_fd_sc_hd__or2_4 c453(
.A(net220),
.B(net396),
.X(out46)
);

sky130_fd_sc_hd__o21ba_2 c454(
.A1(net95),
.A2(net388),
.B1_N(out19),
.X(net400)
);

sky130_fd_sc_hd__nand2b_1 c455(
.A_N(net391),
.B(net651),
.Y(net401)
);

sky130_fd_sc_hd__nor2_1 c456(
.A(net400),
.B(net95),
.Y(out27)
);

sky130_fd_sc_hd__dfrbp_1 c457(
.D(net273),
.RESET_B(out19),
.CLK(clk),
.Q(net402)
);

sky130_fd_sc_hd__nor2_1 c458(
.A(net399),
.B(net401),
.Y(net403)
);

sky130_fd_sc_hd__o21ba_2 c459(
.A1(net403),
.A2(net382),
.B1_N(net395),
.X(net404)
);

sky130_fd_sc_hd__mux4_2 c460(
.A0(net398),
.A1(net265),
.A2(net386),
.A3(net220),
.S0(out11),
.S1(net388),
.X(out37)
);

sky130_fd_sc_hd__nor2_2 c461(
.A(net404),
.B(out37),
.Y(net405)
);

sky130_fd_sc_hd__and2b_4 c462(
.A_N(net99),
.B(out41),
.X(net406)
);

sky130_fd_sc_hd__or2b_4 c463(
.A(net38),
.B_N(out4),
.X(net407)
);

sky130_fd_sc_hd__o21bai_2 c464(
.A1(out32),
.A2(out41),
.B1_N(net645),
.Y(net408)
);

sky130_fd_sc_hd__clkbuf_4 c465(
.A(net665),
.X(net409)
);

sky130_fd_sc_hd__nor2_1 c466(
.A(net369),
.B(net406),
.Y(net410)
);

sky130_fd_sc_hd__inv_6 c467(
.A(net665),
.Y(net411)
);

sky130_fd_sc_hd__sdfbbn_1 c468(
.D(net302),
.RESET_B(net369),
.SCD(out37),
.SCE(net395),
.SET_B(net408),
.CLK_N(clk),
.Q(net412)
);

sky130_fd_sc_hd__o21ba_4 c469(
.A1(net104),
.A2(net406),
.B1_N(net339),
.X(out47)
);

sky130_fd_sc_hd__o21ai_2 c470(
.A1(net396),
.A2(out51),
.B1(net209),
.Y(net413)
);

sky130_fd_sc_hd__sdfxtp_1 c471(
.D(net408),
.SCD(net290),
.SCE(net298),
.CLK(clk),
.Q(net414)
);

sky130_fd_sc_hd__mux4_1 c472(
.A0(net411),
.A1(net408),
.A2(net413),
.A3(out51),
.S0(net406),
.S1(out28),
.X(net415)
);

sky130_fd_sc_hd__and2_2 c473(
.A(net412),
.B(net406),
.X(net416)
);

sky130_fd_sc_hd__sdfxtp_2 c474(
.D(net413),
.SCD(net300),
.SCE(net388),
.CLK(clk),
.Q(net417)
);

sky130_fd_sc_hd__o21ai_4 c475(
.A1(net414),
.A2(net408),
.B1(net396),
.Y(net418)
);

sky130_fd_sc_hd__a21oi_2 c476(
.A1(net416),
.A2(net408),
.B1(net410),
.Y(net419)
);

sky130_fd_sc_hd__o21ai_4 c477(
.A1(net406),
.A2(net417),
.B1(net652),
.Y(out38)
);

sky130_fd_sc_hd__o41a_4 c478(
.A1(net409),
.A2(net406),
.A3(net417),
.A4(out31),
.B1(out28),
.X(net420)
);

sky130_fd_sc_hd__or2b_4 c479(
.A(net402),
.B_N(net419),
.X(net421)
);

sky130_fd_sc_hd__mux4_1 c480(
.A0(net390),
.A1(net418),
.A2(net410),
.A3(net421),
.S0(net413),
.S1(net414),
.X(net422)
);

sky130_fd_sc_hd__mux4_2 c481(
.A0(net417),
.A1(net421),
.A2(net408),
.A3(net298),
.S0(net406),
.S1(net653),
.X(net423)
);

sky130_fd_sc_hd__o31ai_2 c482(
.A1(net410),
.A2(net421),
.A3(net339),
.B1(net654),
.Y(net424)
);

sky130_fd_sc_hd__o31ai_2 c494(
.A1(net296),
.A2(net307),
.A3(out45),
.B1(net318),
.Y(net425)
);

sky130_fd_sc_hd__sdfsbp_1 c495(
.D(net298),
.SCD(net209),
.SCE(net104),
.SET_B(net72),
.CLK(clk),
.Q(out33)
);

sky130_fd_sc_hd__o41a_1 c496(
.A1(net186),
.A2(net311),
.A3(net79),
.A4(net194),
.B1(net304),
.X(out50)
);

sky130_fd_sc_hd__sdfbbn_2 c497(
.D(net309),
.RESET_B(net304),
.SCD(net267),
.SCE(out51),
.SET_B(net298),
.CLK_N(clk),
.Q(net426)
);

sky130_fd_sc_hd__o31ai_4 c498(
.A1(net300),
.A2(out43),
.A3(net307),
.B1(net72),
.Y(out14)
);

sky130_fd_sc_hd__mux4_1 c499(
.A0(net118),
.A1(net318),
.A2(net46),
.A3(out32),
.S0(out43),
.S1(out31),
.X(out13)
);

sky130_fd_sc_hd__sdfbbp_1 c500(
.D(net267),
.RESET_B(net194),
.SCD(net321),
.SCE(out11),
.SET_B(out44),
.CLK(clk),
.Q(out48)
);

sky130_fd_sc_hd__sdfbbn_1 c501(
.D(net426),
.RESET_B(net322),
.SCD(out44),
.SCE(out50),
.SET_B(net420),
.CLK_N(clk),
.Q(out49)
);

sky130_fd_sc_hd__sdfsbp_2 c502(
.D(net425),
.SCD(net186),
.SCE(net72),
.SET_B(out50),
.CLK(clk),
.Q(out42)
);

sky130_fd_sc_hd__sdfbbn_2 c503(
.D(net46),
.RESET_B(net420),
.SCD(out41),
.SCE(net299),
.SET_B(out4),
.CLK_N(clk),
.Q(out2)
);

sky130_fd_sc_hd__buf_2 c504(
.A(in3),
.X(net427)
);

sky130_fd_sc_hd__nor2b_4 c505(
.A(net87),
.B_N(out39),
.Y(net428)
);

sky130_fd_sc_hd__buf_8 c506(
.A(net212),
.X(net429)
);

sky130_fd_sc_hd__nand2b_2 c507(
.A_N(in9),
.B(net87),
.Y(net430)
);

sky130_fd_sc_hd__or2b_4 c508(
.A(net85),
.B_N(net93),
.X(net431)
);

sky130_fd_sc_hd__and2b_4 c509(
.A_N(net430),
.B(net76),
.X(net432)
);

sky130_fd_sc_hd__nor2b_1 c510(
.A(net328),
.B_N(net327),
.Y(net433)
);

sky130_fd_sc_hd__and2_2 c511(
.A(net427),
.B(net433),
.X(net434)
);

sky130_fd_sc_hd__nand2_1 c512(
.A(net429),
.B(net328),
.Y(net435)
);

sky130_fd_sc_hd__nor2_4 c513(
.A(net198),
.B(net431),
.Y(net436)
);

sky130_fd_sc_hd__nand2_4 c514(
.A(net76),
.B(net335),
.Y(net437)
);

sky130_fd_sc_hd__and2b_1 c515(
.A_N(net329),
.B(net88),
.X(net438)
);

sky130_fd_sc_hd__nor2b_4 c516(
.A(net435),
.B_N(net431),
.Y(net439)
);

sky130_fd_sc_hd__and2b_2 c517(
.A_N(net437),
.B(net433),
.X(net440)
);

sky130_fd_sc_hd__dfrbp_2 c518(
.D(net429),
.RESET_B(net440),
.CLK(clk),
.Q(net441)
);

sky130_fd_sc_hd__nand2b_1 c519(
.A_N(net325),
.B(net437),
.Y(net442)
);

sky130_fd_sc_hd__nand2b_4 c520(
.A_N(net435),
.B(net433),
.Y(net443)
);

sky130_fd_sc_hd__nor2b_1 c521(
.A(net436),
.B_N(net212),
.Y(net444)
);

sky130_fd_sc_hd__dfrtn_1 c522(
.D(net434),
.RESET_B(net439),
.CLK_N(clk),
.Q(net445)
);

sky130_fd_sc_hd__or2b_1 c523(
.A(net442),
.B_N(net444),
.X(net446)
);

sky130_fd_sc_hd__or2b_4 c524(
.A(net444),
.B_N(net436),
.X(net447)
);

sky130_fd_sc_hd__and2b_2 c525(
.A_N(in3),
.B(net343),
.X(net448)
);

sky130_fd_sc_hd__o31a_4 c526(
.A1(in40),
.A2(net431),
.A3(net360),
.B1(net326),
.X(net449)
);

sky130_fd_sc_hd__and2b_2 c527(
.A_N(net111),
.B(net337),
.X(net450)
);

sky130_fd_sc_hd__dfrtp_1 c528(
.D(net216),
.RESET_B(net439),
.CLK(clk),
.Q(net451)
);

sky130_fd_sc_hd__nor2_2 c529(
.A(net450),
.B(net451),
.Y(net452)
);

sky130_fd_sc_hd__dfrtp_2 c530(
.D(net443),
.RESET_B(net445),
.CLK(clk),
.Q(net453)
);

sky130_fd_sc_hd__nand2b_2 c531(
.A_N(net326),
.B(net359),
.Y(net454)
);

sky130_fd_sc_hd__dfrtp_4 c532(
.D(net453),
.RESET_B(net428),
.CLK(clk),
.Q(net455)
);

sky130_fd_sc_hd__sdfxtp_4 c533(
.D(net428),
.SCD(net443),
.SCE(net344),
.CLK(clk),
.Q(net456)
);

sky130_fd_sc_hd__or2_4 c534(
.A(net441),
.B(net456),
.X(net457)
);

sky130_fd_sc_hd__or2_2 c535(
.A(net451),
.B(net344),
.X(net458)
);

sky130_fd_sc_hd__dfsbp_1 c536(
.D(net452),
.SET_B(net455),
.CLK(clk),
.Q(net459)
);

sky130_fd_sc_hd__o31ai_2 c537(
.A1(net449),
.A2(net455),
.A3(net344),
.B1(net444),
.Y(net460)
);

sky130_fd_sc_hd__a21oi_4 c538(
.A1(net232),
.A2(net354),
.B1(net449),
.Y(net461)
);

sky130_fd_sc_hd__o21ai_4 c539(
.A1(net431),
.A2(net74),
.B1(in6),
.Y(net462)
);

sky130_fd_sc_hd__a21o_1 c540(
.A1(net354),
.A2(net460),
.B1(net458),
.X(net463)
);

sky130_fd_sc_hd__o21a_1 c541(
.A1(net337),
.A2(net209),
.B1(in40),
.X(net464)
);

sky130_fd_sc_hd__nor2b_2 c542(
.A(net454),
.B_N(net457),
.Y(net465)
);

sky130_fd_sc_hd__and2_0 c543(
.A(net459),
.B(net464),
.X(out26)
);

sky130_fd_sc_hd__mux4_1 c544(
.A0(net432),
.A1(net456),
.A2(net461),
.A3(net352),
.S0(out26),
.S1(net433),
.X(net466)
);

sky130_fd_sc_hd__sdfbbp_1 c545(
.D(net448),
.RESET_B(net343),
.SCD(out26),
.SCE(net359),
.SET_B(net344),
.CLK(clk),
.Q(net468),
.Q_N(net467)
);

sky130_fd_sc_hd__nor2_4 c546(
.A(in6),
.B(net384),
.Y(net469)
);

sky130_fd_sc_hd__or2b_1 c547(
.A(net124),
.B_N(net444),
.X(net470)
);

sky130_fd_sc_hd__and2b_2 c548(
.A_N(net122),
.B(net242),
.X(net471)
);

sky130_fd_sc_hd__and2_0 c549(
.A(net242),
.B(net470),
.X(net472)
);

sky130_fd_sc_hd__dfsbp_2 c550(
.D(net469),
.SET_B(out26),
.CLK(clk),
.Q(net474),
.Q_N(net473)
);

sky130_fd_sc_hd__nor2_1 c551(
.A(net103),
.B(net472),
.Y(net475)
);

sky130_fd_sc_hd__nor2_2 c552(
.A(net343),
.B(net458),
.Y(net476)
);

sky130_fd_sc_hd__a21boi_1 c553(
.A1(net476),
.A2(net127),
.B1_N(net371),
.Y(net477)
);

sky130_fd_sc_hd__nand2_4 c554(
.A(net361),
.B(in6),
.Y(net478)
);

sky130_fd_sc_hd__a21oi_4 c555(
.A1(net355),
.A2(net474),
.B1(net458),
.Y(net479)
);

sky130_fd_sc_hd__and2b_2 c556(
.A_N(net465),
.B(net363),
.X(net480)
);

sky130_fd_sc_hd__mux4_4 c557(
.A0(net332),
.A1(net477),
.A2(net377),
.A3(out26),
.S0(net479),
.S1(net343),
.X(net481)
);

sky130_fd_sc_hd__dfstp_1 c558(
.D(net475),
.SET_B(net127),
.CLK(clk),
.Q(net482)
);

sky130_fd_sc_hd__dfbbn_1 c559(
.D(net479),
.RESET_B(net252),
.SET_B(net471),
.CLK_N(clk),
.Q(net483)
);

sky130_fd_sc_hd__nor2b_2 c560(
.A(net367),
.B_N(net474),
.Y(net484)
);

sky130_fd_sc_hd__sdfstp_1 c561(
.D(net372),
.SCD(net381),
.SCE(net384),
.SET_B(out26),
.CLK(clk),
.Q(net485)
);

sky130_fd_sc_hd__o31ai_4 c562(
.A1(net371),
.A2(net367),
.A3(net485),
.B1(net473),
.Y(net486)
);

sky130_fd_sc_hd__dfstp_2 c563(
.D(net378),
.SET_B(net485),
.CLK(clk),
.Q(net487)
);

sky130_fd_sc_hd__nor2b_4 c564(
.A(net485),
.B_N(net487),
.Y(net488)
);

sky130_fd_sc_hd__o41a_4 c565(
.A1(net480),
.A2(net486),
.A3(net444),
.A4(net487),
.B1(net465),
.X(net489)
);

sky130_fd_sc_hd__mux4_1 c566(
.A0(net471),
.A1(net489),
.A2(net343),
.A3(net132),
.S0(net486),
.S1(net656),
.X(net490)
);

sky130_fd_sc_hd__mux2_8 c567(
.A0(net28),
.A1(net93),
.S(net381),
.X(net491)
);

sky130_fd_sc_hd__dfstp_4 c568(
.D(net491),
.SET_B(out26),
.CLK(clk),
.Q(net492)
);

sky130_fd_sc_hd__dfbbn_2 c569(
.D(in23),
.RESET_B(net252),
.SET_B(net492),
.CLK_N(clk),
.Q(net493)
);

sky130_fd_sc_hd__dfbbp_1 c570(
.D(net440),
.RESET_B(net458),
.SET_B(net491),
.CLK(clk),
.Q(net495),
.Q_N(net494)
);

sky130_fd_sc_hd__and2_1 c571(
.A(net478),
.B(net492),
.X(net496)
);

sky130_fd_sc_hd__a21boi_4 c572(
.A1(net389),
.A2(net491),
.B1_N(net392),
.Y(net497)
);

sky130_fd_sc_hd__sdfxbp_1 c573(
.D(net375),
.SCD(net493),
.SCE(net492),
.CLK(clk),
.Q(net498)
);

sky130_fd_sc_hd__o21ba_2 c574(
.A1(net492),
.A2(net339),
.B1_N(net389),
.X(net499)
);

sky130_fd_sc_hd__mux4_2 c575(
.A0(net496),
.A1(net24),
.A2(net491),
.A3(net388),
.S0(out19),
.S1(net494),
.X(net500)
);

sky130_fd_sc_hd__dlrbn_1 c576(
.D(net381),
.RESET_B(net405),
.GATE_N(clk),
.Q(out5),
.Q_N(net501)
);

sky130_fd_sc_hd__dlrbn_2 c577(
.D(net497),
.RESET_B(net499),
.GATE_N(clk),
.Q(net503),
.Q_N(net502)
);

sky130_fd_sc_hd__o21ai_0 c578(
.A1(net498),
.A2(out29),
.B1(net501),
.Y(net504)
);

sky130_fd_sc_hd__or2b_1 c579(
.A(net359),
.B_N(net502),
.X(net505)
);

sky130_fd_sc_hd__and2b_4 c580(
.A_N(net505),
.B(out5),
.X(net506)
);

sky130_fd_sc_hd__o31ai_1 c581(
.A1(net135),
.A2(net506),
.A3(net381),
.B1(net501),
.Y(net507)
);

sky130_fd_sc_hd__or2b_1 c582(
.A(net339),
.B_N(net503),
.X(net508)
);

sky130_fd_sc_hd__nand2b_2 c583(
.A_N(net504),
.B(net506),
.Y(net509)
);

sky130_fd_sc_hd__nand2b_1 c584(
.A_N(net507),
.B(net470),
.Y(net510)
);

sky130_fd_sc_hd__sdfxbp_2 c585(
.D(net508),
.SCD(net510),
.SCE(net458),
.CLK(clk),
.Q(net511)
);

sky130_fd_sc_hd__or2_1 c586(
.A(net383),
.B(net509),
.X(net512)
);

sky130_fd_sc_hd__mux4_2 c587(
.A0(net512),
.A1(net511),
.A2(net507),
.A3(net509),
.S0(net382),
.S1(net494),
.X(net513)
);

sky130_fd_sc_hd__o21ai_1 c588(
.A1(net503),
.A2(net363),
.B1(in13),
.Y(net514)
);

sky130_fd_sc_hd__or2_4 c589(
.A(net407),
.B(net509),
.X(net515)
);

sky130_fd_sc_hd__o21ba_1 c590(
.A1(net487),
.A2(net506),
.B1_N(out30),
.X(net516)
);

sky130_fd_sc_hd__dlygate4sd3_1 c591(
.A(net664),
.X(net517)
);

sky130_fd_sc_hd__a21o_4 c592(
.A1(net155),
.A2(net421),
.B1(out32),
.X(net518)
);

sky130_fd_sc_hd__o21ai_4 c593(
.A1(net141),
.A2(out5),
.B1(out29),
.Y(net519)
);

sky130_fd_sc_hd__a21bo_4 c594(
.A1(net482),
.A2(net339),
.B1_N(net458),
.X(net520)
);

sky130_fd_sc_hd__a21o_2 c595(
.A1(net392),
.A2(out37),
.B1(net509),
.X(net521)
);

sky130_fd_sc_hd__clkbuf_1 c596(
.A(net664),
.X(out25)
);

sky130_fd_sc_hd__mux4_2 c597(
.A0(net166),
.A1(net517),
.A2(net506),
.A3(out25),
.S0(out37),
.S1(net407),
.X(net522)
);

sky130_fd_sc_hd__sdfstp_2 c598(
.D(net520),
.SCD(net474),
.SCE(net513),
.SET_B(out25),
.CLK(clk),
.Q(net523)
);

sky130_fd_sc_hd__mux4_4 c599(
.A0(net519),
.A1(net171),
.A2(in18),
.A3(out25),
.S0(net473),
.S1(net517),
.X(net524)
);

sky130_fd_sc_hd__o31a_1 c600(
.A1(net281),
.A2(net388),
.A3(out38),
.B1(net657),
.X(net525)
);

sky130_fd_sc_hd__o21ba_4 c601(
.A1(net446),
.A2(net474),
.B1_N(net658),
.X(net526)
);

sky130_fd_sc_hd__sdfxtp_1 c602(
.D(net252),
.SCD(net525),
.SCE(in18),
.CLK(clk),
.Q(net527)
);

sky130_fd_sc_hd__sdfxtp_2 c603(
.D(net518),
.SCD(out25),
.SCE(net509),
.CLK(clk),
.Q(net528)
);

sky130_fd_sc_hd__sdfstp_4 c604(
.D(net527),
.SCD(net526),
.SCE(out26),
.SET_B(out11),
.CLK(clk),
.Q(out36)
);

sky130_fd_sc_hd__sdfxtp_4 c605(
.D(net363),
.SCD(net513),
.SCE(net204),
.CLK(clk),
.Q(net529)
);

sky130_fd_sc_hd__sdfbbn_1 c606(
.D(net500),
.RESET_B(out25),
.SCD(net513),
.SCE(net526),
.SET_B(net171),
.CLK_N(clk),
.Q(net530)
);

sky130_fd_sc_hd__a21boi_2 c607(
.A1(net528),
.A2(net458),
.B1_N(out29),
.Y(net531)
);

sky130_fd_sc_hd__a21o_2 c608(
.A1(net495),
.A2(net529),
.B1(net531),
.X(net532)
);

sky130_fd_sc_hd__and2b_4 c630(
.A_N(net324),
.B(out39),
.X(net533)
);

sky130_fd_sc_hd__and2_0 c631(
.A(net438),
.B(net445),
.X(net534)
);

sky130_fd_sc_hd__clkbuf_1 c632(
.A(net637),
.X(net535)
);

sky130_fd_sc_hd__inv_2 c633(
.A(net637),
.Y(net536)
);

sky130_fd_sc_hd__dlrbp_1 c634(
.D(net439),
.RESET_B(net204),
.GATE(clk),
.Q(net538),
.Q_N(net537)
);

sky130_fd_sc_hd__nand2_4 c635(
.A(in5),
.B(net534),
.Y(net539)
);

sky130_fd_sc_hd__and2b_4 c636(
.A_N(in18),
.B(net445),
.X(net540)
);

sky130_fd_sc_hd__nor2_1 c637(
.A(in20),
.B(net537),
.Y(net541)
);

sky130_fd_sc_hd__dlrbp_2 c638(
.D(net88),
.RESET_B(net434),
.GATE(clk),
.Q(net543),
.Q_N(net542)
);

sky130_fd_sc_hd__nand2b_2 c639(
.A_N(net534),
.B(out39),
.Y(net544)
);

sky130_fd_sc_hd__or2_2 c640(
.A(net535),
.B(net542),
.X(net545)
);

sky130_fd_sc_hd__nand2b_1 c641(
.A_N(net543),
.B(in20),
.Y(net546)
);

sky130_fd_sc_hd__dlrtn_1 c642(
.D(net334),
.RESET_B(net534),
.GATE_N(clk),
.Q(net547)
);

sky130_fd_sc_hd__dlrtn_2 c643(
.D(net338),
.RESET_B(net209),
.GATE_N(clk),
.Q(net548)
);

sky130_fd_sc_hd__nor2b_1 c644(
.A(net548),
.B_N(net541),
.Y(net549)
);

sky130_fd_sc_hd__and2_2 c645(
.A(net547),
.B(net539),
.X(net550)
);

sky130_fd_sc_hd__dlrtn_4 c646(
.D(net544),
.RESET_B(net545),
.GATE_N(clk),
.Q(net551)
);

sky130_fd_sc_hd__o21ba_2 c647(
.A1(net550),
.A2(net551),
.B1_N(net537),
.X(net552)
);

sky130_fd_sc_hd__dlrtp_1 c648(
.D(net552),
.RESET_B(net538),
.GATE(clk),
.Q(net553)
);

sky130_fd_sc_hd__a21o_1 c649(
.A1(net553),
.A2(net438),
.B1(net548),
.X(net554)
);

sky130_fd_sc_hd__dfbbn_1 c650(
.D(net534),
.RESET_B(net554),
.SET_B(net552),
.CLK_N(clk),
.Q(net556),
.Q_N(net555)
);

sky130_fd_sc_hd__and2_4 c651(
.A(net461),
.B(in14),
.X(net557)
);

sky130_fd_sc_hd__and2_2 c652(
.A(net113),
.B(net538),
.X(net558)
);

sky130_fd_sc_hd__dlrtp_2 c653(
.D(net540),
.RESET_B(net557),
.GATE(clk),
.Q(net559)
);

sky130_fd_sc_hd__o41a_4 c654(
.A1(net457),
.A2(out4),
.A3(net558),
.A4(net468),
.B1(net541),
.X(net560)
);

sky130_fd_sc_hd__nand2_4 c655(
.A(net558),
.B(net93),
.Y(net561)
);

sky130_fd_sc_hd__mux4_1 c656(
.A0(net352),
.A1(net468),
.A2(net555),
.A3(in5),
.S0(net558),
.S1(net557),
.X(net562)
);

sky130_fd_sc_hd__or2_2 c657(
.A(net238),
.B(net540),
.X(net563)
);

sky130_fd_sc_hd__dlrtp_4 c658(
.D(net462),
.RESET_B(net557),
.GATE(clk),
.Q(net564)
);

sky130_fd_sc_hd__edfxbp_1 c659(
.D(net557),
.DE(net546),
.CLK(clk),
.Q(net565)
);

sky130_fd_sc_hd__or2b_4 c660(
.A(net463),
.B_N(net558),
.X(net566)
);

sky130_fd_sc_hd__and2_2 c661(
.A(net565),
.B(net462),
.X(net567)
);

sky130_fd_sc_hd__mux4_2 c662(
.A0(net561),
.A1(net209),
.A2(out39),
.A3(net557),
.S0(net563),
.S1(net238),
.X(net568)
);

sky130_fd_sc_hd__or2_4 c663(
.A(net468),
.B(net564),
.X(net569)
);

sky130_fd_sc_hd__and2b_1 c664(
.A_N(net566),
.B(net564),
.X(net570)
);

sky130_fd_sc_hd__and2_0 c665(
.A(net556),
.B(net655),
.X(net571)
);

sky130_fd_sc_hd__and2_4 c666(
.A(net560),
.B(net571),
.X(net572)
);

sky130_fd_sc_hd__mux4_1 c667(
.A0(net347),
.A1(out39),
.A2(net557),
.A3(out23),
.S0(net570),
.S1(net549),
.X(net573)
);

sky130_fd_sc_hd__o21ai_4 c668(
.A1(net570),
.A2(net467),
.B1(net659),
.Y(net574)
);

sky130_fd_sc_hd__sdfbbn_2 c669(
.D(net439),
.RESET_B(net558),
.SCD(net467),
.SCE(net464),
.SET_B(net661),
.CLK_N(clk),
.Q(net575)
);

sky130_fd_sc_hd__mux4_1 c670(
.A0(net464),
.A1(net558),
.A2(net541),
.A3(net536),
.S0(net433),
.S1(net660),
.X(net576)
);

sky130_fd_sc_hd__edfxtp_1 c671(
.D(net576),
.DE(net575),
.CLK(clk),
.Q(net577)
);

sky130_fd_sc_hd__nor2_4 c672(
.A(net445),
.B(net549),
.Y(net578)
);

sky130_fd_sc_hd__or2b_4 c673(
.A(net569),
.B_N(net537),
.X(out15)
);

sky130_fd_sc_hd__nand2b_2 c674(
.A_N(net572),
.B(out39),
.Y(net579)
);

sky130_fd_sc_hd__and2b_1 c675(
.A_N(net559),
.B(net570),
.X(net580)
);

sky130_fd_sc_hd__o41a_4 c676(
.A1(net538),
.A2(net489),
.A3(out39),
.A4(net577),
.B1(net563),
.X(net581)
);

sky130_fd_sc_hd__dfbbn_2 c677(
.D(net377),
.RESET_B(net581),
.SET_B(in14),
.CLK_N(clk),
.Q(net582)
);

sky130_fd_sc_hd__dfbbp_1 c678(
.D(net483),
.RESET_B(net581),
.SET_B(net577),
.CLK(clk),
.Q(net584),
.Q_N(net583)
);

sky130_fd_sc_hd__a21oi_1 c679(
.A1(net132),
.A2(net551),
.B1(net541),
.Y(net585)
);

sky130_fd_sc_hd__sedfxbp_1 c680(
.D(net582),
.DE(net581),
.SCD(net489),
.SCE(net377),
.CLK(clk),
.Q(net586)
);

sky130_fd_sc_hd__sdfxbp_1 c681(
.D(net578),
.SCD(net464),
.SCE(net581),
.CLK(clk),
.Q(net587)
);

sky130_fd_sc_hd__inv_1 c682(
.A(net642),
.Y(net588)
);

sky130_fd_sc_hd__inv_12 c683(
.A(net641),
.Y(net589)
);

sky130_fd_sc_hd__o21ai_0 c684(
.A1(net545),
.A2(net588),
.B1(net577),
.Y(net590)
);

sky130_fd_sc_hd__sdfxbp_2 c685(
.D(net580),
.SCD(net590),
.SCE(net588),
.CLK(clk),
.Q(net592),
.Q_N(net591)
);

sky130_fd_sc_hd__sdfxtp_1 c686(
.D(net585),
.SCD(net592),
.SCE(net580),
.CLK(clk),
.Q(net593)
);

sky130_fd_sc_hd__o41a_4 c687(
.A1(net127),
.A2(net593),
.A3(out15),
.A4(net590),
.B1(net584),
.X(net594)
);

sky130_fd_sc_hd__o41a_4 c688(
.A1(net567),
.A2(net589),
.A3(net445),
.A4(net577),
.B1(net488),
.X(net595)
);

sky130_fd_sc_hd__o21bai_4 c689(
.A1(net551),
.A2(net589),
.B1_N(net595),
.Y(out12)
);

sky130_fd_sc_hd__o31a_1 c690(
.A1(net484),
.A2(net595),
.A3(out12),
.B1(net594),
.X(net596)
);

sky130_fd_sc_hd__o41a_2 c691(
.A1(net384),
.A2(net595),
.A3(net464),
.A4(net591),
.B1(net563),
.X(net597)
);

sky130_fd_sc_hd__mux2_4 c692(
.A0(net594),
.A1(out12),
.S(net595),
.X(net598)
);

sky130_fd_sc_hd__buf_6 c693(
.A(net663),
.X(out7)
);

sky130_fd_sc_hd__buf_12 c694(
.A(net663),
.X(net599)
);

sky130_fd_sc_hd__sdfxtp_2 c695(
.D(net564),
.SCD(net277),
.SCE(out19),
.CLK(clk),
.Q(out1)
);

sky130_fd_sc_hd__o21bai_2 c696(
.A1(net563),
.A2(net145),
.B1_N(out23),
.Y(net600)
);

sky130_fd_sc_hd__o21a_2 c697(
.A1(net433),
.A2(out6),
.B1(in41),
.X(net601)
);

sky130_fd_sc_hd__sdfxtp_4 c698(
.D(net601),
.SCD(out4),
.SCE(net495),
.CLK(clk),
.Q(net602)
);

sky130_fd_sc_hd__mux4_2 c699(
.A0(net570),
.A1(net592),
.A2(net433),
.A3(out15),
.S0(net494),
.S1(net577),
.X(net603)
);

sky130_fd_sc_hd__a21o_4 c700(
.A1(net536),
.A2(in14),
.B1(net570),
.X(net604)
);

sky130_fd_sc_hd__dfbbn_1 c701(
.D(net79),
.RESET_B(net604),
.SET_B(net564),
.CLK_N(clk),
.Q(net605)
);

sky130_fd_sc_hd__or2b_2 c702(
.A(net464),
.B_N(net596),
.X(net606)
);

sky130_fd_sc_hd__dfbbn_2 c703(
.D(net606),
.RESET_B(net495),
.SET_B(out5),
.CLK_N(clk),
.Q(net608),
.Q_N(net607)
);

sky130_fd_sc_hd__dfbbp_1 c704(
.D(net277),
.RESET_B(net577),
.SET_B(net601),
.CLK(clk),
.Q(net610),
.Q_N(net609)
);

sky130_fd_sc_hd__and2_0 c705(
.A(net610),
.B(net495),
.X(net611)
);

sky130_fd_sc_hd__a21o_4 c706(
.A1(net587),
.A2(net21),
.B1(net607),
.X(net612)
);

sky130_fd_sc_hd__mux4_4 c707(
.A0(net600),
.A1(net145),
.A2(net609),
.A3(net591),
.S0(net501),
.S1(net570),
.X(net613)
);

sky130_fd_sc_hd__mux2_2 c708(
.A0(net24),
.A1(net605),
.S(net564),
.X(net614)
);

sky130_fd_sc_hd__a21o_2 c709(
.A1(net541),
.A2(net599),
.B1(net209),
.X(out17)
);

sky130_fd_sc_hd__mux2_2 c710(
.A0(net612),
.A1(net611),
.S(net464),
.X(net615)
);

sky130_fd_sc_hd__mux4_1 c711(
.A0(net613),
.A1(net574),
.A2(net546),
.A3(net489),
.S0(net564),
.S1(net596),
.X(net616)
);

sky130_fd_sc_hd__a21oi_2 c712(
.A1(net614),
.A2(net584),
.B1(net662),
.Y(net617)
);

sky130_fd_sc_hd__sdfxbp_1 c713(
.D(net608),
.SCD(in13),
.SCE(net581),
.CLK(clk),
.Q(net618)
);

sky130_fd_sc_hd__a21bo_1 c714(
.A1(net516),
.A2(net93),
.B1_N(out19),
.X(net619)
);

sky130_fd_sc_hd__inv_16 c715(
.A(net635),
.Y(out16)
);

sky130_fd_sc_hd__sedfxbp_2 c716(
.D(net549),
.DE(net615),
.SCD(net489),
.SCE(net546),
.CLK(clk),
.Q(net620)
);

sky130_fd_sc_hd__o41a_4 c717(
.A1(net209),
.A2(net530),
.A3(net598),
.A4(net93),
.B1(out4),
.X(net621)
);

sky130_fd_sc_hd__o31a_1 c718(
.A1(net488),
.A2(net523),
.A3(net388),
.B1(net204),
.X(net622)
);

sky130_fd_sc_hd__mux2_8 c719(
.A0(net602),
.A1(net489),
.S(out23),
.X(net623)
);

sky130_fd_sc_hd__o21a_4 c720(
.A1(net447),
.A2(net619),
.B1(out12),
.X(net624)
);

sky130_fd_sc_hd__clkinv_1 c721(
.A(net635),
.Y(net625)
);

sky130_fd_sc_hd__sedfxtp_1 c722(
.D(net93),
.DE(net590),
.SCD(net447),
.SCE(net424),
.CLK(clk),
.Q(net626)
);

sky130_fd_sc_hd__o31a_2 c723(
.A1(net620),
.A2(net626),
.A3(net488),
.B1(net657),
.X(net627)
);

sky130_fd_sc_hd__sdfxbp_2 c724(
.D(net623),
.SCD(net624),
.SCE(net204),
.CLK(clk),
.Q(net628)
);

sky130_fd_sc_hd__o21a_2 c725(
.A1(net546),
.A2(net598),
.B1(net626),
.X(net629)
);

sky130_fd_sc_hd__o21a_2 c726(
.A1(net628),
.A2(net618),
.B1(in41),
.X(net630)
);

sky130_fd_sc_hd__o41a_2 c727(
.A1(net627),
.A2(net625),
.A3(out6),
.A4(net447),
.B1(net501),
.X(net631)
);

sky130_fd_sc_hd__mux4_4 c728(
.A0(net586),
.A1(net631),
.A2(net629),
.A3(net626),
.S0(out1),
.S1(net657),
.X(out18)
);

sky130_fd_sc_hd__sdfxtp_1 c729(
.D(net581),
.SCD(net621),
.SCE(out15),
.CLK(clk),
.Q(out10)
);

sky130_fd_sc_hd__a21boi_4 c730(
.A1(net629),
.A2(net622),
.B1_N(out8),
.Y(net632)
);

sky130_fd_sc_hd__o21ai_1 c731(
.A1(in41),
.A2(net532),
.B1(out8),
.Y(net633)
);

sky130_fd_sc_hd__o31ai_2 c732(
.A1(net630),
.A2(net515),
.A3(out8),
.B1(net626),
.Y(net634)
);

sky130_fd_sc_hd__o31ai_4 c733(
.A1(net633),
.A2(net617),
.A3(net447),
.B1(net629),
.Y(out3)
);

sky130_fd_sc_hd__sdfxtp_2 c734(
.D(net634),
.SCD(net632),
.SCE(net629),
.CLK(clk)
);

sky130_fd_sc_hd__sedfxtp_2 merge755(
.D(net539),
.DE(net603),
.SCD(net424),
.SCE(net388),
.CLK(clk),
.Q(net635)
);

sky130_fd_sc_hd__mux4_4 merge756(
.A0(net117),
.A1(net597),
.A2(net464),
.A3(net583),
.S0(net494),
.S1(net581),
.X(net636)
);

sky130_fd_sc_hd__sedfxtp_4 merge757(
.D(net74),
.DE(net439),
.SCD(net533),
.SCE(net433),
.CLK(clk),
.Q(net637)
);

sky130_fd_sc_hd__sdfrbp_1 merge758(
.D(net152),
.RESET_B(net40),
.SCD(net44),
.SCE(net157),
.CLK(clk),
.Q(net639),
.Q_N(net638)
);

sky130_fd_sc_hd__mux4_2 merge759(
.A0(net514),
.A1(net473),
.A2(net500),
.A3(net521),
.S0(out32),
.S1(net166),
.X(net640)
);

sky130_fd_sc_hd__sdfrbp_2 merge760(
.D(net579),
.RESET_B(net132),
.SCD(net490),
.SCE(net580),
.CLK(clk),
.Q(net642),
.Q_N(net641)
);

sky130_fd_sc_hd__mux4_1 merge761(
.A0(net114),
.A1(net302),
.A2(net141),
.A3(net290),
.S0(net171),
.S1(out6),
.X(net643)
);

sky130_fd_sc_hd__dfxbp_1 s762(
.D(net173),
.CLK(clk),
.Q(net645),
.Q_N(net644)
);

sky130_fd_sc_hd__dfxbp_2 s763(
.D(net187),
.CLK(clk),
.Q(net646)
);

sky130_fd_sc_hd__dfxtp_1 s764(
.D(net193),
.CLK(clk),
.Q(net647)
);

sky130_fd_sc_hd__dfxtp_2 s765(
.D(net253),
.CLK(clk),
.Q(net648)
);

sky130_fd_sc_hd__dfxtp_4 s766(
.D(net257),
.CLK(clk),
.Q(net649)
);

sky130_fd_sc_hd__dlclkp_1 s767(
.GATE(net268),
.CLK(clk),
.GCLK(net650)
);

sky130_fd_sc_hd__dlclkp_2 s768(
.GATE(net278),
.CLK(clk),
.GCLK(net651)
);

sky130_fd_sc_hd__dlclkp_4 s769(
.GATE(net415),
.CLK(clk),
.GCLK(net652)
);

sky130_fd_sc_hd__dlxbn_1 s770(
.D(net422),
.GATE_N(clk),
.Q(net653)
);

sky130_fd_sc_hd__dlxbn_2 s771(
.D(net423),
.GATE_N(clk),
.Q(net654)
);

sky130_fd_sc_hd__dlxbp_1 s772(
.D(net466),
.GATE(clk),
.Q(net655)
);

sky130_fd_sc_hd__dlxtn_1 s773(
.D(net481),
.GATE_N(clk),
.Q(net656)
);

sky130_fd_sc_hd__dlxtn_2 s774(
.D(net522),
.GATE_N(clk),
.Q(net657)
);

sky130_fd_sc_hd__dlxtn_4 s775(
.D(net524),
.GATE_N(clk),
.Q(net658)
);

sky130_fd_sc_hd__dlxtp_1 s776(
.D(net562),
.GATE(clk),
.Q(net659)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s777(
.D(net568),
.SLEEP_B(clk),
.Q(net660)
);

sky130_fd_sc_hd__dfxbp_1 s778(
.D(net573),
.CLK(clk),
.Q(net661)
);

sky130_fd_sc_hd__dfxbp_2 s779(
.D(net616),
.CLK(clk),
.Q(net662)
);

sky130_fd_sc_hd__dfxtp_1 s780(
.D(net636),
.CLK(clk),
.Q(net663)
);

sky130_fd_sc_hd__dfxtp_2 s781(
.D(net640),
.CLK(clk),
.Q(net664)
);

sky130_fd_sc_hd__dfxtp_4 s782(
.D(net643),
.CLK(clk),
.Q(net665)
);


endmodule
