module netlist_1 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input in52,
	input in53,
	input in54,
	input in55,
	input in56,
	input in57,
	input in58,
	input in59,
	input in60,
	input in61,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51,
	output out52,
	output out53,
	output out54,
	output out55,
	output out56,
	output out57,
	output out58,
	output out59,
	output out60,
	output out61
);


wire clk;
wire net731;
wire net730;
wire net729;
wire net728;
wire net726;
wire net725;
wire net724;
wire net722;
wire net720;
wire net719;
wire net717;
wire net716;
wire net715;
wire net714;
wire net712;
wire net711;
wire net708;
wire net706;
wire net705;
wire net704;
wire net703;
wire net701;
wire net699;
wire out3;
wire net698;
wire net697;
wire net696;
wire net695;
wire out11;
wire net694;
wire net693;
wire net692;
wire net690;
wire out20;
wire net687;
wire net686;
wire net685;
wire net684;
wire net683;
wire net680;
wire net671;
wire net669;
wire net668;
wire net370;
wire net667;
wire net664;
wire net659;
wire in6;
wire net656;
wire out53;
wire out58;
wire out49;
wire net462;
wire out7;
wire net652;
wire net622;
wire net651;
wire out17;
wire out23;
wire net304;
wire net645;
wire net641;
wire out38;
wire net637;
wire net632;
wire net665;
wire net631;
wire net629;
wire net74;
wire net628;
wire net3;
wire net627;
wire net447;
wire net626;
wire net624;
wire net506;
wire net623;
wire net620;
wire in49;
wire net619;
wire net46;
wire net615;
wire net347;
wire net100;
wire net288;
wire net614;
wire net165;
wire net613;
wire net20;
wire net612;
wire net638;
wire net428;
wire net610;
wire out25;
wire net608;
wire net1;
wire net424;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire net601;
wire net596;
wire net592;
wire net588;
wire net587;
wire in4;
wire net583;
wire net707;
wire net582;
wire net158;
wire net584;
wire net581;
wire net336;
wire net579;
wire net577;
wire net576;
wire out2;
wire net570;
wire net209;
wire net569;
wire in41;
wire net567;
wire in30;
wire net566;
wire net565;
wire net39;
wire net562;
wire net559;
wire net556;
wire net647;
wire net555;
wire net159;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire in55;
wire net550;
wire net710;
wire net544;
wire net539;
wire net534;
wire net532;
wire net271;
wire net530;
wire net617;
wire net306;
wire net537;
wire net369;
wire net528;
wire net525;
wire net523;
wire net520;
wire net519;
wire net516;
wire net672;
wire net514;
wire net78;
wire net508;
wire net721;
wire net504;
wire net679;
wire out57;
wire net503;
wire net573;
wire net224;
wire net499;
wire net674;
wire net496;
wire net495;
wire net494;
wire net179;
wire in39;
wire net453;
wire net493;
wire net472;
wire net492;
wire net479;
wire net491;
wire net295;
wire net490;
wire net489;
wire net487;
wire net486;
wire net478;
wire net474;
wire net473;
wire net468;
wire net540;
wire net202;
wire net465;
wire net469;
wire net471;
wire net461;
wire net546;
wire net460;
wire net454;
wire out13;
wire net648;
wire net452;
wire net449;
wire net448;
wire net498;
wire net700;
wire net446;
wire net691;
wire net88;
wire net444;
wire in59;
wire net110;
wire net442;
wire net609;
wire net440;
wire net128;
wire net439;
wire net147;
wire out21;
wire net438;
wire net433;
wire net432;
wire out41;
wire net419;
wire net431;
wire net430;
wire net618;
wire net429;
wire net427;
wire net426;
wire net673;
wire net425;
wire net423;
wire net183;
wire net531;
wire net421;
wire net52;
wire net170;
wire net420;
wire net450;
wire net418;
wire net415;
wire net414;
wire net276;
wire net413;
wire net330;
wire net252;
wire net412;
wire net411;
wire net517;
wire net677;
wire net410;
wire net409;
wire net407;
wire out19;
wire net406;
wire net662;
wire net405;
wire net607;
wire net526;
wire net404;
wire net29;
wire net403;
wire net383;
wire net663;
wire net402;
wire net106;
wire net572;
wire net401;
wire net399;
wire net398;
wire out46;
wire net476;
wire net396;
wire net172;
wire net395;
wire net391;
wire net443;
wire net557;
wire net345;
wire net527;
wire net488;
wire net390;
wire net441;
wire out15;
wire out5;
wire net646;
wire net389;
wire net513;
wire net501;
wire out14;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net131;
wire net184;
wire net380;
wire net379;
wire net260;
wire net616;
wire net378;
wire net543;
wire net38;
wire net377;
wire net376;
wire net625;
wire net373;
wire net598;
wire net374;
wire out37;
wire net676;
wire net372;
wire net371;
wire net368;
wire net367;
wire net366;
wire net365;
wire net364;
wire net363;
wire net360;
wire net660;
wire out28;
wire net359;
wire net397;
wire net357;
wire net356;
wire net510;
wire net355;
wire net521;
wire net353;
wire net590;
wire net507;
wire net351;
wire net350;
wire out30;
wire net547;
wire net511;
wire net451;
wire net13;
wire net343;
wire net89;
wire net666;
wire net340;
wire net339;
wire net337;
wire net458;
wire net538;
wire net244;
wire net334;
wire net333;
wire net332;
wire net331;
wire net328;
wire net327;
wire net119;
wire net325;
wire net324;
wire net321;
wire net535;
wire net320;
wire net542;
wire net139;
wire net318;
wire out9;
wire net335;
wire net315;
wire net313;
wire net505;
wire net199;
wire out27;
wire net294;
wire net319;
wire net312;
wire net309;
wire net308;
wire net417;
wire net302;
wire net298;
wire net296;
wire in24;
wire net358;
wire net127;
wire net293;
wire in56;
wire net134;
wire out48;
wire net305;
wire net594;
wire out39;
wire net292;
wire net230;
wire out22;
wire net500;
wire net445;
wire net303;
wire net291;
wire net201;
wire net422;
wire net289;
wire net595;
wire net384;
wire net482;
wire in25;
wire net286;
wire net153;
wire out61;
wire net589;
wire net278;
wire net274;
wire net643;
wire net273;
wire net142;
wire out10;
wire net272;
wire net114;
wire net270;
wire in17;
wire net267;
wire net644;
wire net266;
wire net459;
wire net463;
wire net0;
wire net297;
wire net408;
wire net475;
wire net280;
wire net102;
wire net151;
wire net275;
wire net264;
wire net657;
wire net591;
wire net196;
wire net262;
wire net217;
wire net261;
wire net21;
wire net257;
wire net689;
wire net44;
wire net117;
wire net62;
wire net109;
wire net254;
wire net203;
wire net253;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire in26;
wire net661;
wire net194;
wire net241;
wire out42;
wire net238;
wire net234;
wire net232;
wire out12;
wire net226;
wire out32;
wire net568;
wire net375;
wire net223;
wire net524;
wire net575;
wire net382;
wire net548;
wire net259;
wire net222;
wire net31;
wire net219;
wire net578;
wire net210;
wire net326;
wire net213;
wire net208;
wire out16;
wire net188;
wire net207;
wire net649;
wire net205;
wire net678;
wire net633;
wire net122;
wire net197;
wire net483;
wire net193;
wire net192;
wire net190;
wire net630;
wire in20;
wire net189;
wire net246;
wire net186;
wire net152;
wire net126;
wire net113;
wire net284;
wire net655;
wire net563;
wire net464;
wire net549;
wire net182;
wire in29;
wire net240;
wire net416;
wire net41;
wire net104;
wire net8;
wire out33;
wire net310;
wire net180;
wire out40;
wire net258;
wire net176;
wire net342;
wire net17;
wire net437;
wire out44;
wire in35;
wire out24;
wire net580;
wire net133;
wire net175;
wire net80;
wire net173;
wire out52;
wire net195;
wire in37;
wire net518;
wire net381;
wire net218;
wire net300;
wire net169;
wire net485;
wire net344;
wire net168;
wire out6;
wire net167;
wire net509;
wire net58;
wire net221;
wire net166;
wire net269;
wire net97;
wire net434;
wire net204;
wire net200;
wire net621;
wire net162;
wire net316;
wire out31;
wire out60;
wire net497;
wire out45;
wire net161;
wire net285;
wire net160;
wire net636;
wire net311;
wire net150;
wire net149;
wire net111;
wire net124;
wire net242;
wire net290;
wire net227;
wire out47;
wire net148;
wire net178;
wire net239;
wire net144;
wire net322;
wire net688;
wire net299;
wire net143;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net561;
wire out29;
wire net137;
wire net136;
wire net456;
wire net135;
wire net255;
wire net157;
wire net177;
wire net349;
wire out51;
wire net130;
wire in12;
wire net103;
wire net481;
wire net120;
wire net455;
wire net65;
wire net129;
wire net392;
wire out0;
wire net164;
wire net642;
wire net268;
wire in7;
wire net400;
wire net82;
wire net2;
wire net123;
wire net282;
wire net71;
wire net229;
wire in43;
wire net108;
wire net107;
wire out26;
wire net99;
wire net348;
wire net341;
wire in52;
wire net96;
wire net225;
wire net250;
wire net466;
wire net118;
wire net94;
wire net90;
wire net174;
wire net277;
wire net639;
wire net81;
wire in10;
wire net156;
wire net361;
wire net115;
wire net670;
wire in18;
wire net27;
wire net34;
wire net585;
wire net79;
wire net75;
wire net231;
wire net329;
wire net212;
wire net653;
wire in5;
wire net14;
wire net77;
wire net600;
wire net236;
wire net76;
wire in42;
wire net354;
wire in38;
wire net198;
wire net467;
wire net101;
wire net9;
wire net571;
wire net73;
wire net60;
wire net564;
wire net154;
wire net84;
wire in46;
wire net85;
wire net72;
wire net116;
wire net69;
wire net67;
wire in31;
wire net98;
wire net522;
wire net436;
wire net541;
wire net323;
wire net15;
wire net279;
wire net64;
wire net63;
wire net681;
wire net61;
wire net512;
wire net18;
wire out34;
wire net682;
wire net237;
wire net59;
wire net228;
wire net675;
wire net56;
wire net55;
wire net214;
wire net53;
wire in48;
wire net640;
wire net50;
wire net597;
wire out55;
wire net185;
wire net155;
wire net338;
wire net599;
wire net112;
wire net650;
wire net560;
wire net45;
wire net502;
wire net235;
wire net49;
wire in50;
wire net215;
wire net484;
wire net30;
wire out36;
wire in8;
wire net346;
wire net4;
wire net43;
wire net248;
wire net477;
wire out56;
wire net187;
wire in13;
wire net586;
wire net533;
wire net32;
wire net125;
wire net19;
wire in15;
wire net727;
wire net163;
wire in19;
wire net702;
wire net70;
wire net48;
wire net28;
wire net92;
wire net713;
wire net25;
wire in0;
wire net709;
wire net24;
wire net470;
wire in33;
wire net33;
wire net233;
wire net121;
wire net40;
wire in60;
wire net435;
wire net301;
wire net23;
wire net26;
wire net16;
wire net558;
wire in1;
wire net265;
wire net22;
wire net263;
wire net457;
wire out50;
wire net6;
wire net5;
wire net206;
wire in58;
wire in61;
wire net171;
wire in23;
wire out4;
wire net42;
wire net91;
wire in57;
wire net281;
wire net54;
wire in54;
wire out43;
wire in53;
wire net138;
wire net145;
wire net211;
wire net132;
wire in34;
wire net593;
wire in45;
wire net393;
wire net256;
wire net87;
wire net181;
wire net7;
wire out1;
wire out54;
wire net574;
wire net216;
wire out59;
wire in28;
wire in44;
wire in32;
wire net47;
wire net12;
wire in27;
wire in9;
wire net654;
wire net723;
wire net611;
wire net515;
wire net362;
wire in16;
wire net191;
wire net35;
wire net220;
wire in22;
wire net68;
wire in14;
wire net529;
wire in21;
wire net57;
wire net480;
wire net86;
wire net317;
wire in51;
wire net93;
wire in47;
wire in2;
wire net718;
wire net658;
wire net105;
wire in11;
wire net51;
wire in36;
wire net536;
wire net37;
wire net36;
wire net95;
wire net146;
wire net251;
wire net11;
wire net352;
wire net307;
wire net394;
wire net314;
wire in3;
sky130_fd_sc_hd__mux4_1 c62(
.A0(in44),
.A1(in53),
.A2(in57),
.A3(in6),
.S0(in37),
.S1(in54),
.X(net0)
);

sky130_fd_sc_hd__nor2b_2 c63(
.A(in48),
.B_N(net3),
.Y(net1)
);

sky130_fd_sc_hd__nand2_2 c64(
.A(in47),
.B(in54),
.Y(net2)
);

sky130_fd_sc_hd__or3_4 c65(
.A(in38),
.B(in61),
.C(in3),
.X(net3)
);

sky130_fd_sc_hd__and2b_2 c66(
.A_N(in4),
.B(net3),
.X(net4)
);

sky130_fd_sc_hd__and2_0 c67(
.A(in49),
.B(net2),
.X(net5)
);

sky130_fd_sc_hd__nor2b_2 c68(
.A(net2),
.B_N(net4),
.Y(net6)
);

sky130_fd_sc_hd__nor2_4 c69(
.A(net3),
.B(in61),
.Y(net7)
);

sky130_fd_sc_hd__nand2b_1 c70(
.A_N(net5),
.B(net2),
.Y(net8)
);

sky130_fd_sc_hd__or4bb_2 c71(
.A(in60),
.B(net8),
.C_N(net3),
.D_N(net1),
.X(net9)
);

sky130_fd_sc_hd__nand2b_2 c72(
.A_N(net9),
.B(net4),
.Y(net10)
);

sky130_fd_sc_hd__nor2_1 c73(
.A(net5),
.B(in45),
.Y(net11)
);

sky130_fd_sc_hd__nor2_2 c74(
.A(net1),
.B(net9),
.Y(net12)
);

sky130_fd_sc_hd__nand2_4 c75(
.A(net4),
.B(net3),
.Y(net13)
);

sky130_fd_sc_hd__or2_4 c76(
.A(in37),
.B(net0),
.X(net14)
);

sky130_fd_sc_hd__and2_2 c77(
.A(in26),
.B(net13),
.X(net15)
);

sky130_fd_sc_hd__o2111ai_2 c78(
.A1(net11),
.A2(in32),
.B1(in40),
.C1(net13),
.D1(net15),
.Y(net16)
);

sky130_fd_sc_hd__nand2_1 c79(
.A(net8),
.B(net14),
.Y(net17)
);

sky130_fd_sc_hd__and2_4 c80(
.A(in0),
.B(net16),
.X(net18)
);

sky130_fd_sc_hd__o2111ai_2 c81(
.A1(in45),
.A2(net7),
.B1(net18),
.C1(net15),
.D1(net14),
.Y(net19)
);

sky130_fd_sc_hd__or4bb_4 c82(
.A(net17),
.B(net15),
.C_N(net5),
.D_N(net14),
.X(net20)
);

sky130_fd_sc_hd__mux4_1 c83(
.A0(net16),
.A1(net17),
.A2(net20),
.A3(net14),
.S0(net13),
.S1(net19),
.X(net21)
);

sky130_fd_sc_hd__or2b_1 c84(
.A(net16),
.B_N(net14),
.X(net22)
);

sky130_fd_sc_hd__and2b_4 c85(
.A_N(net2),
.B(net4),
.X(net23)
);

sky130_fd_sc_hd__or2_4 c86(
.A(in52),
.B(net16),
.X(net24)
);

sky130_fd_sc_hd__nand2b_2 c87(
.A_N(in25),
.B(in11),
.Y(net25)
);

sky130_fd_sc_hd__or4bb_1 c88(
.A(net24),
.B(net14),
.C_N(net12),
.D_N(net8),
.X(net26)
);

sky130_fd_sc_hd__and2_0 c89(
.A(net4),
.B(net25),
.X(net27)
);

sky130_fd_sc_hd__and2_0 c90(
.A(net6),
.B(net25),
.X(net28)
);

sky130_fd_sc_hd__nand2_4 c91(
.A(in53),
.B(net23),
.Y(net29)
);

sky130_fd_sc_hd__or2_2 c92(
.A(in32),
.B(in50),
.X(net30)
);

sky130_fd_sc_hd__or2_1 c93(
.A(net22),
.B(net25),
.X(net31)
);

sky130_fd_sc_hd__nand2_2 c94(
.A(net25),
.B(net28),
.Y(net32)
);

sky130_fd_sc_hd__and2_1 c95(
.A(net29),
.B(net25),
.X(net33)
);

sky130_fd_sc_hd__o2111a_2 c96(
.A1(net27),
.A2(net33),
.B1(net4),
.C1(in21),
.D1(net28),
.X(net34)
);

sky130_fd_sc_hd__mux4_4 c97(
.A0(net31),
.A1(net13),
.A2(net6),
.A3(net24),
.S0(net25),
.S1(net30),
.X(out51)
);

sky130_fd_sc_hd__or2b_4 c98(
.A(net7),
.B_N(net31),
.X(net35)
);

sky130_fd_sc_hd__nor2_2 c99(
.A(net28),
.B(net33),
.Y(net36)
);

sky130_fd_sc_hd__mux4_4 c100(
.A0(net23),
.A1(net33),
.A2(net34),
.A3(net16),
.S0(net35),
.S1(in22),
.X(net37)
);

sky130_fd_sc_hd__nor2_1 c101(
.A(in15),
.B(net33),
.Y(net38)
);

sky130_fd_sc_hd__mux4_1 c102(
.A0(in57),
.A1(net37),
.A2(in22),
.A3(net38),
.S0(out51),
.S1(net13),
.X(net39)
);

sky130_fd_sc_hd__nor3b_2 c103(
.A(net37),
.B(net39),
.C_N(out51),
.Y(out56)
);

sky130_fd_sc_hd__mux4_1 c104(
.A0(net39),
.A1(net35),
.A2(net33),
.A3(out56),
.S0(net34),
.S1(net38),
.X(net40)
);

sky130_fd_sc_hd__or2_4 c105(
.A(net12),
.B(out56),
.X(net41)
);

sky130_fd_sc_hd__and2_2 c106(
.A(in44),
.B(out51),
.X(net42)
);

sky130_fd_sc_hd__or2b_2 c107(
.A(net41),
.B_N(in32),
.X(net43)
);

sky130_fd_sc_hd__or2_2 c108(
.A(in33),
.B(net32),
.X(net44)
);

sky130_fd_sc_hd__nand2_1 c109(
.A(net11),
.B(out56),
.Y(net45)
);

sky130_fd_sc_hd__and2b_1 c110(
.A_N(net43),
.B(out56),
.X(net46)
);

sky130_fd_sc_hd__nand2_1 c111(
.A(net33),
.B(net44),
.Y(net47)
);

sky130_fd_sc_hd__nand2b_2 c112(
.A_N(in34),
.B(net33),
.Y(net48)
);

sky130_fd_sc_hd__and2_2 c113(
.A(in40),
.B(in50),
.X(net49)
);

sky130_fd_sc_hd__nor2_1 c114(
.A(in32),
.B(net47),
.Y(net50)
);

sky130_fd_sc_hd__nand2b_1 c115(
.A_N(net50),
.B(net48),
.Y(net51)
);

sky130_fd_sc_hd__or4bb_2 c116(
.A(net51),
.B(net8),
.C_N(net49),
.D_N(net32),
.X(net52)
);

sky130_fd_sc_hd__nand2b_1 c117(
.A_N(net49),
.B(net52),
.Y(net53)
);

sky130_fd_sc_hd__and2_2 c118(
.A(net46),
.B(out56),
.X(net54)
);

sky130_fd_sc_hd__or2_1 c119(
.A(net47),
.B(net52),
.X(net55)
);

sky130_fd_sc_hd__mux4_4 c120(
.A0(net54),
.A1(net55),
.A2(net49),
.A3(net50),
.S0(net43),
.S1(net44),
.X(net56)
);

sky130_fd_sc_hd__or2_2 c121(
.A(net48),
.B(net49),
.X(net57)
);

sky130_fd_sc_hd__a2111o_1 c122(
.A1(net44),
.A2(net47),
.B1(net55),
.C1(net43),
.D1(net8),
.X(net58)
);

sky130_fd_sc_hd__or4bb_1 c123(
.A(net57),
.B(net55),
.C_N(net58),
.D_N(net46),
.X(net59)
);

sky130_fd_sc_hd__mux4_4 c124(
.A0(net59),
.A1(net52),
.A2(net57),
.A3(net54),
.S0(out51),
.S1(in17),
.X(net60)
);

sky130_fd_sc_hd__dfrbp_1 c125(
.D(net53),
.RESET_B(net59),
.CLK(clk),
.Q(net62),
.Q_N(net61)
);

sky130_fd_sc_hd__nand2b_2 c126(
.A_N(in7),
.B(in1),
.Y(net63)
);

sky130_fd_sc_hd__and3_2 c127(
.A(in18),
.B(in3),
.C(in11),
.X(net64)
);

sky130_fd_sc_hd__nor3b_4 c128(
.A(in20),
.B(in6),
.C_N(in11),
.Y(net65)
);

sky130_fd_sc_hd__mux4_2 c129(
.A0(in15),
.A1(in1),
.A2(in19),
.A3(in11),
.S0(net63),
.S1(in17),
.X(net66)
);

sky130_fd_sc_hd__and3_4 c130(
.A(net65),
.B(in16),
.C(in17),
.X(net67)
);

sky130_fd_sc_hd__and3b_2 c131(
.A_N(net63),
.B(in17),
.C(in12),
.X(net68)
);

sky130_fd_sc_hd__and3_4 c132(
.A(net66),
.B(in18),
.C(in10),
.X(net69)
);

sky130_fd_sc_hd__nor3b_2 c133(
.A(net66),
.B(net69),
.C_N(in12),
.Y(net70)
);

sky130_fd_sc_hd__a2111oi_0 c134(
.A1(net63),
.A2(in8),
.B1(in13),
.C1(in6),
.D1(in17),
.Y(net71)
);

sky130_fd_sc_hd__nor3_4 c135(
.A(in7),
.B(net71),
.C(net64),
.Y(net72)
);

sky130_fd_sc_hd__o2111a_1 c136(
.A1(net66),
.A2(in8),
.B1(net72),
.C1(net63),
.D1(net68),
.X(net73)
);

sky130_fd_sc_hd__nand3_4 c137(
.A(net68),
.B(in7),
.C(net63),
.Y(net74)
);

sky130_fd_sc_hd__or2b_4 c138(
.A(net67),
.B_N(in20),
.X(net75)
);

sky130_fd_sc_hd__or4bb_2 c139(
.A(net73),
.B(net67),
.C_N(in17),
.D_N(in12),
.X(net76)
);

sky130_fd_sc_hd__nor3_2 c140(
.A(net70),
.B(in18),
.C(in11),
.Y(net77)
);

sky130_fd_sc_hd__nand3b_2 c141(
.A_N(net74),
.B(in3),
.C(net76),
.Y(net78)
);

sky130_fd_sc_hd__mux4_1 c142(
.A0(net69),
.A1(net75),
.A2(net78),
.A3(net68),
.S0(net66),
.S1(net67),
.X(net79)
);

sky130_fd_sc_hd__nor3_1 c143(
.A(net79),
.B(net67),
.C(net77),
.Y(net80)
);

sky130_fd_sc_hd__a2111oi_2 c144(
.A1(net76),
.A2(net78),
.B1(in0),
.C1(net75),
.D1(in17),
.Y(net81)
);

sky130_fd_sc_hd__mux4_1 c145(
.A0(net80),
.A1(net81),
.A2(net75),
.A3(net74),
.S0(net66),
.S1(net77),
.X(net82)
);

sky130_fd_sc_hd__mux4_4 c146(
.A0(net66),
.A1(net82),
.A2(net76),
.A3(net65),
.S0(net74),
.S1(in17),
.X(net83)
);

sky130_fd_sc_hd__or4bb_4 c147(
.A(in31),
.B(in16),
.C_N(in33),
.D_N(net76),
.X(net84)
);

sky130_fd_sc_hd__nand3b_1 c148(
.A_N(net64),
.B(in12),
.C(net83),
.Y(net85)
);

sky130_fd_sc_hd__or3b_1 c149(
.A(net84),
.B(in6),
.C_N(in17),
.X(net86)
);

sky130_fd_sc_hd__and3_2 c150(
.A(net70),
.B(in25),
.C(net63),
.X(net87)
);

sky130_fd_sc_hd__and2b_4 c151(
.A_N(net87),
.B(net78),
.X(net88)
);

sky130_fd_sc_hd__or4bb_1 c152(
.A(in24),
.B(in25),
.C_N(in36),
.D_N(net78),
.X(net89)
);

sky130_fd_sc_hd__and2_1 c153(
.A(net82),
.B(in9),
.X(net90)
);

sky130_fd_sc_hd__mux4_2 c154(
.A0(net90),
.A1(net72),
.A2(in14),
.A3(net86),
.S0(in25),
.S1(in41),
.X(net91)
);

sky130_fd_sc_hd__nor2_1 c155(
.A(in35),
.B(net90),
.Y(net92)
);

sky130_fd_sc_hd__or2_4 c156(
.A(net83),
.B(net90),
.X(net93)
);

sky130_fd_sc_hd__nand3b_2 c157(
.A_N(net93),
.B(net84),
.C(net85),
.Y(net94)
);

sky130_fd_sc_hd__nand3b_1 c158(
.A_N(in28),
.B(net92),
.C(net91),
.Y(net95)
);

sky130_fd_sc_hd__a2111oi_2 c159(
.A1(in12),
.A2(net89),
.B1(net90),
.C1(net94),
.D1(net81),
.Y(net96)
);

sky130_fd_sc_hd__nor2_2 c160(
.A(in13),
.B(net92),
.Y(net97)
);

sky130_fd_sc_hd__o2111a_2 c161(
.A1(net95),
.A2(net97),
.B1(net78),
.C1(in28),
.D1(net81),
.X(net98)
);

sky130_fd_sc_hd__and3_1 c162(
.A(net98),
.B(in12),
.C(net95),
.X(net99)
);

sky130_fd_sc_hd__or4bb_2 c163(
.A(net99),
.B(net98),
.C_N(in17),
.D_N(net88),
.X(net100)
);

sky130_fd_sc_hd__sdfrbp_1 c164(
.D(net96),
.RESET_B(in29),
.SCD(net100),
.SCE(net90),
.CLK(clk),
.Q(net102),
.Q_N(net101)
);

sky130_fd_sc_hd__mux4_2 c165(
.A0(net92),
.A1(net100),
.A2(net98),
.A3(net97),
.S0(net91),
.S1(net70),
.X(net103)
);

sky130_fd_sc_hd__mux4_2 c166(
.A0(net94),
.A1(net89),
.A2(net91),
.A3(net90),
.S0(net98),
.S1(net639),
.X(net104)
);

sky130_fd_sc_hd__mux4_2 c167(
.A0(net94),
.A1(net100),
.A2(net95),
.A3(net96),
.S0(net74),
.S1(net639),
.X(net105)
);

sky130_fd_sc_hd__nand3_2 c168(
.A(net75),
.B(in43),
.C(net101),
.Y(net106)
);

sky130_fd_sc_hd__nor2b_2 c169(
.A(net79),
.B_N(in6),
.Y(net107)
);

sky130_fd_sc_hd__or3_2 c170(
.A(net104),
.B(net106),
.C(net78),
.X(net108)
);

sky130_fd_sc_hd__sdfrbp_2 c171(
.D(in43),
.RESET_B(net108),
.SCD(net75),
.SCE(in51),
.CLK(clk),
.Q(net110),
.Q_N(net109)
);

sky130_fd_sc_hd__nor3b_4 c172(
.A(net102),
.B(net107),
.C_N(in56),
.Y(net111)
);

sky130_fd_sc_hd__and2b_2 c173(
.A_N(net106),
.B(net107),
.X(net112)
);

sky130_fd_sc_hd__and2_1 c174(
.A(net78),
.B(net111),
.X(net113)
);

sky130_fd_sc_hd__and2_0 c175(
.A(net111),
.B(in55),
.X(net114)
);

sky130_fd_sc_hd__nand2b_2 c176(
.A_N(net65),
.B(net113),
.Y(net115)
);

sky130_fd_sc_hd__mux4_1 c177(
.A0(net110),
.A1(net106),
.A2(net75),
.A3(net112),
.S0(net79),
.S1(net84),
.X(net116)
);

sky130_fd_sc_hd__dfbbn_1 c178(
.D(net108),
.RESET_B(net112),
.SET_B(net114),
.CLK_N(clk),
.Q(net118),
.Q_N(net117)
);

sky130_fd_sc_hd__nand3b_1 c179(
.A_N(in1),
.B(in27),
.C(net102),
.Y(net119)
);

sky130_fd_sc_hd__mux4_2 c180(
.A0(net116),
.A1(net96),
.A2(net91),
.A3(net117),
.S0(net109),
.S1(net114),
.X(net120)
);

sky130_fd_sc_hd__or3b_4 c181(
.A(net120),
.B(net106),
.C_N(net115),
.X(net121)
);

sky130_fd_sc_hd__sdfbbn_1 c182(
.D(net113),
.RESET_B(net121),
.SCD(net120),
.SCE(net112),
.SET_B(in51),
.CLK_N(clk),
.Q(net123),
.Q_N(net122)
);

sky130_fd_sc_hd__sdfbbn_2 c183(
.D(net118),
.RESET_B(net120),
.SCD(net114),
.SCE(net116),
.SET_B(net121),
.CLK_N(clk),
.Q(net125),
.Q_N(net124)
);

sky130_fd_sc_hd__mux4_4 c184(
.A0(net115),
.A1(net120),
.A2(net111),
.A3(net96),
.S0(in55),
.S1(net121),
.X(net126)
);

sky130_fd_sc_hd__dfbbn_2 c185(
.D(net121),
.RESET_B(net124),
.SET_B(net641),
.CLK_N(clk),
.Q(net128),
.Q_N(net127)
);

sky130_fd_sc_hd__mux4_2 c186(
.A0(in42),
.A1(net121),
.A2(net112),
.A3(net127),
.S0(net124),
.S1(net641),
.X(net129)
);

sky130_fd_sc_hd__mux4_4 c187(
.A0(net107),
.A1(net114),
.A2(in55),
.A3(net0),
.S0(net641),
.S1(net642),
.X(net130)
);

sky130_fd_sc_hd__mux4_1 c188(
.A0(net130),
.A1(net108),
.A2(net128),
.A3(net122),
.S0(net120),
.S1(net641),
.X(net131)
);

sky130_fd_sc_hd__nor2b_2 c189(
.A(net10),
.B_N(net19),
.Y(net132)
);

sky130_fd_sc_hd__sdfrtn_1 c190(
.D(in25),
.RESET_B(net10),
.SCD(net121),
.SCE(net642),
.CLK_N(clk),
.Q(net133)
);

sky130_fd_sc_hd__a2111oi_2 c191(
.A1(in46),
.A2(net0),
.B1(net133),
.C1(in17),
.D1(in0),
.Y(net134)
);

sky130_fd_sc_hd__nand2b_4 c192(
.A_N(net15),
.B(net20),
.Y(net135)
);

sky130_fd_sc_hd__nand3b_1 c193(
.A_N(net19),
.B(net125),
.C(net135),
.Y(net136)
);

sky130_fd_sc_hd__nor2b_2 c194(
.A(net134),
.B_N(net88),
.Y(net137)
);

sky130_fd_sc_hd__o2111ai_4 c195(
.A1(net0),
.A2(net21),
.B1(net137),
.C1(net74),
.D1(net135),
.Y(net138)
);

sky130_fd_sc_hd__and3b_2 c196(
.A_N(in3),
.B(net19),
.C(net10),
.X(net139)
);

sky130_fd_sc_hd__nor3_4 c197(
.A(in55),
.B(net134),
.C(net139),
.Y(net140)
);

sky130_fd_sc_hd__a2111o_1 c198(
.A1(net133),
.A2(net74),
.B1(in46),
.C1(net135),
.D1(net139),
.X(net141)
);

sky130_fd_sc_hd__or4bb_1 c199(
.A(net135),
.B(net88),
.C_N(net139),
.D_N(net642),
.X(net142)
);

sky130_fd_sc_hd__or4bb_4 c200(
.A(net135),
.B(net139),
.C_N(net142),
.D_N(net642),
.X(net143)
);

sky130_fd_sc_hd__o2111a_2 c201(
.A1(net139),
.A2(net135),
.B1(net15),
.C1(net141),
.D1(net142),
.X(net144)
);

sky130_fd_sc_hd__mux4_1 c202(
.A0(net132),
.A1(net21),
.A2(net135),
.A3(net138),
.S0(net143),
.S1(net142),
.X(net145)
);

sky130_fd_sc_hd__or4bb_2 c203(
.A(net143),
.B(net139),
.C_N(net124),
.D_N(net142),
.X(net146)
);

sky130_fd_sc_hd__nand3_4 c204(
.A(net136),
.B(net15),
.C(net142),
.Y(net147)
);

sky130_fd_sc_hd__mux4_2 c205(
.A0(net138),
.A1(net135),
.A2(net144),
.A3(net145),
.S0(net14),
.S1(net127),
.X(net148)
);

sky130_fd_sc_hd__mux4_4 c206(
.A0(net141),
.A1(net140),
.A2(net125),
.A3(net146),
.S0(net139),
.S1(net142),
.X(out47)
);

sky130_fd_sc_hd__and3_2 c207(
.A(net21),
.B(net139),
.C(net142),
.X(net149)
);

sky130_fd_sc_hd__mux4_2 c208(
.A0(net144),
.A1(net149),
.A2(net132),
.A3(net135),
.S0(net139),
.S1(net145),
.X(out55)
);

sky130_fd_sc_hd__mux4_4 c209(
.A0(net149),
.A1(net145),
.A2(net138),
.A3(net135),
.S0(net142),
.S1(net139),
.X(net150)
);

sky130_fd_sc_hd__mux4_2 c210(
.A0(net31),
.A1(net34),
.A2(net14),
.A3(net148),
.S0(net146),
.S1(net25),
.X(out29)
);

sky130_fd_sc_hd__nand2b_2 c211(
.A_N(net26),
.B(net8),
.Y(net151)
);

sky130_fd_sc_hd__or2b_1 c212(
.A(net140),
.B_N(net137),
.X(net152)
);

sky130_fd_sc_hd__nor2b_4 c213(
.A(net152),
.B_N(net74),
.Y(net153)
);

sky130_fd_sc_hd__nand2b_2 c214(
.A_N(net137),
.B(net97),
.Y(net154)
);

sky130_fd_sc_hd__nand3b_1 c215(
.A_N(net148),
.B(net97),
.C(net38),
.Y(net155)
);

sky130_fd_sc_hd__a2111oi_4 c216(
.A1(net81),
.A2(in4),
.B1(net38),
.C1(out56),
.D1(net145),
.Y(net156)
);

sky130_fd_sc_hd__a2111o_1 c217(
.A1(net88),
.A2(net128),
.B1(net137),
.C1(net8),
.D1(net152),
.X(net157)
);

sky130_fd_sc_hd__and3b_2 c218(
.A_N(net25),
.B(net137),
.C(in5),
.X(net158)
);

sky130_fd_sc_hd__and3_2 c219(
.A(net151),
.B(net25),
.C(in54),
.X(net159)
);

sky130_fd_sc_hd__nor3b_1 c220(
.A(net35),
.B(net147),
.C_N(net27),
.Y(net160)
);

sky130_fd_sc_hd__nor2b_2 c221(
.A(net158),
.B_N(net27),
.Y(net161)
);

sky130_fd_sc_hd__or2_1 c222(
.A(net160),
.B(net152),
.X(out31)
);

sky130_fd_sc_hd__nor3_4 c223(
.A(net97),
.B(in4),
.C(in56),
.Y(out60)
);

sky130_fd_sc_hd__and2b_2 c224(
.A_N(net125),
.B(net155),
.X(net162)
);

sky130_fd_sc_hd__mux4_1 c225(
.A0(in4),
.A1(net161),
.A2(in11),
.A3(net38),
.S0(out60),
.S1(net36),
.X(net163)
);

sky130_fd_sc_hd__o2111ai_4 c226(
.A1(net162),
.A2(net13),
.B1(net147),
.C1(net40),
.D1(net31),
.Y(out26)
);

sky130_fd_sc_hd__nand3b_1 c227(
.A_N(net74),
.B(net162),
.C(net160),
.Y(net164)
);

sky130_fd_sc_hd__and2b_1 c228(
.A_N(net153),
.B(net145),
.X(net165)
);

sky130_fd_sc_hd__and3b_2 c229(
.A_N(net165),
.B(net160),
.C(out31),
.X(out42)
);

sky130_fd_sc_hd__mux4_4 c230(
.A0(net30),
.A1(net138),
.A2(net97),
.A3(net165),
.S0(out42),
.S1(net25),
.X(net166)
);

sky130_fd_sc_hd__nor3b_4 c231(
.A(net52),
.B(out60),
.C_N(net43),
.Y(out39)
);

sky130_fd_sc_hd__or3b_1 c232(
.A(net42),
.B(net156),
.C_N(out60),
.X(net167)
);

sky130_fd_sc_hd__nand3b_2 c233(
.A_N(net147),
.B(net138),
.C(net638),
.Y(out6)
);

sky130_fd_sc_hd__nand3_2 c234(
.A(net166),
.B(out47),
.C(out59),
.Y(net168)
);

sky130_fd_sc_hd__o2111a_1 c235(
.A1(net156),
.A2(out39),
.B1(net58),
.C1(net47),
.D1(net8),
.X(net169)
);

sky130_fd_sc_hd__or4bb_1 c236(
.A(net43),
.B(net147),
.C_N(net161),
.D_N(net32),
.X(net170)
);

sky130_fd_sc_hd__a2111oi_2 c237(
.A1(net62),
.A2(net49),
.B1(net58),
.C1(net42),
.D1(net638),
.Y(net171)
);

sky130_fd_sc_hd__and3b_4 c238(
.A_N(net170),
.B(out6),
.C(net52),
.X(net172)
);

sky130_fd_sc_hd__nor3_1 c239(
.A(net32),
.B(net166),
.C(net170),
.Y(out10)
);

sky130_fd_sc_hd__sdfbbp_1 c240(
.D(net63),
.RESET_B(in33),
.SCD(out10),
.SCE(out26),
.SET_B(net161),
.CLK(clk),
.Q(net174),
.Q_N(net173)
);

sky130_fd_sc_hd__sdfbbn_1 c241(
.D(net161),
.RESET_B(out26),
.SCD(out31),
.SCE(out56),
.SET_B(net173),
.CLK_N(clk),
.Q(out24),
.Q_N(net175)
);

sky130_fd_sc_hd__sdfrtp_1 c242(
.D(net174),
.RESET_B(out39),
.SCD(out10),
.SCE(net175),
.CLK(clk),
.Q(out44)
);

sky130_fd_sc_hd__o2111ai_1 c243(
.A1(net55),
.A2(net47),
.B1(net62),
.C1(in54),
.D1(net138),
.Y(net176)
);

sky130_fd_sc_hd__mux4_4 c244(
.A0(net172),
.A1(net169),
.A2(out55),
.A3(net147),
.S0(net42),
.S1(out31),
.X(net177)
);

sky130_fd_sc_hd__a2111o_4 c245(
.A1(in11),
.A2(out24),
.B1(net63),
.C1(net147),
.D1(out38),
.X(out54)
);

sky130_fd_sc_hd__dfbbp_1 c246(
.D(net168),
.RESET_B(out6),
.SET_B(net637),
.CLK(clk),
.Q(out34),
.Q_N(net178)
);

sky130_fd_sc_hd__sdfbbn_2 c247(
.D(net45),
.RESET_B(out34),
.SCD(net175),
.SCE(net61),
.SET_B(net169),
.CLK_N(clk),
.Q(out57),
.Q_N(net179)
);

sky130_fd_sc_hd__or4bb_1 c248(
.A(net167),
.B(out57),
.C_N(net55),
.D_N(net45),
.X(net180)
);

sky130_fd_sc_hd__sdfbbp_1 c249(
.D(net171),
.RESET_B(net43),
.SCD(out57),
.SCE(net178),
.SET_B(net176),
.CLK(clk),
.Q(out33)
);

sky130_fd_sc_hd__sdfrtp_2 c250(
.D(net180),
.RESET_B(out10),
.SCD(net174),
.SCE(net179),
.CLK(clk),
.Q(net181)
);

sky130_fd_sc_hd__and3_4 c251(
.A(net181),
.B(net63),
.C(net179),
.X(net182)
);

sky130_fd_sc_hd__nor2b_2 c252(
.A(in11),
.B_N(net68),
.Y(net183)
);

sky130_fd_sc_hd__or4bb_4 c253(
.A(in8),
.B(net77),
.C_N(in6),
.D_N(net69),
.X(net184)
);

sky130_fd_sc_hd__and2b_1 c254(
.A_N(net183),
.B(net77),
.X(net185)
);

sky130_fd_sc_hd__or2_1 c255(
.A(net67),
.B(in2),
.X(net186)
);

sky130_fd_sc_hd__nor2b_2 c256(
.A(net185),
.B_N(net186),
.Y(net187)
);

sky130_fd_sc_hd__nor2b_4 c257(
.A(in5),
.B_N(net183),
.Y(net188)
);

sky130_fd_sc_hd__or2_2 c258(
.A(net187),
.B(net188),
.X(net189)
);

sky130_fd_sc_hd__o2111ai_4 c259(
.A1(net77),
.A2(net69),
.B1(net71),
.C1(net184),
.D1(net68),
.Y(net190)
);

sky130_fd_sc_hd__or4bb_4 c260(
.A(in19),
.B(net184),
.C_N(net67),
.D_N(in17),
.X(out40)
);

sky130_fd_sc_hd__mux4_4 c261(
.A0(net73),
.A1(net189),
.A2(net187),
.A3(net184),
.S0(net186),
.S1(net188),
.X(net191)
);

sky130_fd_sc_hd__nor3_2 c262(
.A(net183),
.B(net190),
.C(net186),
.Y(net192)
);

sky130_fd_sc_hd__a2111oi_0 c263(
.A1(net186),
.A2(in2),
.B1(net184),
.C1(net191),
.D1(in0),
.Y(net193)
);

sky130_fd_sc_hd__o2111a_2 c264(
.A1(net189),
.A2(net184),
.B1(net193),
.C1(net191),
.D1(net190),
.X(net194)
);

sky130_fd_sc_hd__mux4_1 c265(
.A0(in20),
.A1(in11),
.A2(net77),
.A3(in6),
.S0(net184),
.S1(net187),
.X(net195)
);

sky130_fd_sc_hd__or2_1 c266(
.A(in10),
.B(net194),
.X(net196)
);

sky130_fd_sc_hd__mux4_2 c267(
.A0(net195),
.A1(net194),
.A2(net191),
.A3(in19),
.S0(net189),
.S1(net183),
.X(net197)
);

sky130_fd_sc_hd__or3_2 c268(
.A(out40),
.B(net193),
.C(net188),
.X(net198)
);

sky130_fd_sc_hd__mux4_2 c269(
.A0(net192),
.A1(net187),
.A2(net67),
.A3(out40),
.S0(net195),
.S1(net196),
.X(net199)
);

sky130_fd_sc_hd__and2_4 c270(
.A(net197),
.B(net72),
.X(out1)
);

sky130_fd_sc_hd__mux4_1 c271(
.A0(net193),
.A1(net199),
.A2(net188),
.A3(net196),
.S0(net187),
.S1(net191),
.X(net200)
);

sky130_fd_sc_hd__nor3b_1 c272(
.A(net199),
.B(net186),
.C_N(net197),
.Y(net201)
);

sky130_fd_sc_hd__nor2b_2 c273(
.A(net76),
.B_N(out40),
.Y(net202)
);

sky130_fd_sc_hd__nor2b_2 c274(
.A(net72),
.B_N(net96),
.Y(net203)
);

sky130_fd_sc_hd__and2_2 c275(
.A(in2),
.B(in9),
.X(net204)
);

sky130_fd_sc_hd__dfrbp_2 c276(
.D(in29),
.RESET_B(net100),
.CLK(clk),
.Q(net206),
.Q_N(net205)
);

sky130_fd_sc_hd__nand2b_4 c277(
.A_N(net89),
.B(in14),
.Y(net207)
);

sky130_fd_sc_hd__and2_2 c278(
.A(net204),
.B(net76),
.X(net208)
);

sky130_fd_sc_hd__or2_4 c279(
.A(net207),
.B(net89),
.X(net209)
);

sky130_fd_sc_hd__nand2b_4 c280(
.A_N(in9),
.B(net204),
.Y(net210)
);

sky130_fd_sc_hd__or4bb_2 c281(
.A(net210),
.B(net76),
.C_N(net190),
.D_N(in17),
.X(net211)
);

sky130_fd_sc_hd__a2111o_4 c282(
.A1(net190),
.A2(net209),
.B1(net208),
.C1(in23),
.D1(net640),
.X(net212)
);

sky130_fd_sc_hd__or4bb_2 c283(
.A(net208),
.B(net76),
.C_N(net206),
.D_N(net211),
.X(net213)
);

sky130_fd_sc_hd__or3_2 c284(
.A(net208),
.B(net188),
.C(net205),
.X(net214)
);

sky130_fd_sc_hd__sdfrtp_4 c285(
.D(net211),
.RESET_B(net202),
.SCD(net100),
.SCE(out1),
.CLK(clk),
.Q(net215)
);

sky130_fd_sc_hd__mux4_4 c286(
.A0(net215),
.A1(net204),
.A2(net212),
.A3(net209),
.S0(net100),
.S1(net210),
.X(net216)
);

sky130_fd_sc_hd__and2b_1 c287(
.A_N(net203),
.B(net89),
.X(net217)
);

sky130_fd_sc_hd__sdfbbn_1 c288(
.D(net100),
.RESET_B(net203),
.SCD(net212),
.SCE(net89),
.SET_B(net198),
.CLK_N(clk),
.Q(net219),
.Q_N(net218)
);

sky130_fd_sc_hd__nor2_4 c289(
.A(net219),
.B(net209),
.Y(net220)
);

sky130_fd_sc_hd__mux4_4 c290(
.A0(net214),
.A1(net209),
.A2(net72),
.A3(net202),
.S0(net212),
.S1(net644),
.X(net221)
);

sky130_fd_sc_hd__a2111oi_0 c291(
.A1(net214),
.A2(net219),
.B1(net207),
.C1(net72),
.D1(net191),
.Y(net222)
);

sky130_fd_sc_hd__mux4_2 c292(
.A0(net222),
.A1(net215),
.A2(net72),
.A3(net196),
.S0(net217),
.S1(net645),
.X(net223)
);

sky130_fd_sc_hd__mux4_1 c293(
.A0(net217),
.A1(net214),
.A2(net218),
.A3(net222),
.S0(net215),
.S1(out23),
.X(net224)
);

sky130_fd_sc_hd__nand3b_4 c294(
.A_N(in6),
.B(net119),
.C(net643),
.Y(net225)
);

sky130_fd_sc_hd__nand3b_1 c295(
.A_N(in58),
.B(net122),
.C(net205),
.Y(net226)
);

sky130_fd_sc_hd__nor2_1 c296(
.A(net196),
.B(net647),
.Y(net227)
);

sky130_fd_sc_hd__and2_0 c297(
.A(net119),
.B(net643),
.X(net228)
);

sky130_fd_sc_hd__mux4_2 c298(
.A0(net114),
.A1(net227),
.A2(net228),
.A3(net226),
.S0(in27),
.S1(in17),
.X(net229)
);

sky130_fd_sc_hd__or4bb_2 c299(
.A(in51),
.B(net206),
.C_N(net123),
.D_N(net648),
.X(net230)
);

sky130_fd_sc_hd__or2_2 c300(
.A(in59),
.B(in21),
.X(net231)
);

sky130_fd_sc_hd__nor2b_1 c301(
.A(net91),
.B_N(net227),
.Y(net232)
);

sky130_fd_sc_hd__and3b_4 c302(
.A_N(net231),
.B(net98),
.C(net226),
.X(net233)
);

sky130_fd_sc_hd__nand2_2 c303(
.A(net226),
.B(net114),
.Y(net234)
);

sky130_fd_sc_hd__nand3b_4 c304(
.A_N(net225),
.B(net234),
.C(net215),
.Y(net235)
);

sky130_fd_sc_hd__or3_4 c305(
.A(net235),
.B(net212),
.C(in51),
.X(net236)
);

sky130_fd_sc_hd__nand3b_1 c306(
.A_N(in30),
.B(net234),
.C(net235),
.Y(net237)
);

sky130_fd_sc_hd__nor3b_1 c307(
.A(net229),
.B(net235),
.C_N(net222),
.Y(net238)
);

sky130_fd_sc_hd__nor2_1 c308(
.A(net230),
.B(net127),
.Y(net239)
);

sky130_fd_sc_hd__and2_2 c309(
.A(net236),
.B(net235),
.X(net240)
);

sky130_fd_sc_hd__nand3_4 c310(
.A(net226),
.B(net235),
.C(net233),
.Y(net241)
);

sky130_fd_sc_hd__mux4_4 c311(
.A0(net233),
.A1(net241),
.A2(net119),
.A3(net240),
.S0(net98),
.S1(net236),
.X(net242)
);

sky130_fd_sc_hd__mux4_2 c312(
.A0(net239),
.A1(net235),
.A2(net241),
.A3(net234),
.S0(out40),
.S1(out17),
.X(net243)
);

sky130_fd_sc_hd__sdfsbp_1 c313(
.D(net232),
.SCD(net241),
.SCE(out17),
.SET_B(net649),
.CLK(clk),
.Q(net245),
.Q_N(net244)
);

sky130_fd_sc_hd__mux4_1 c314(
.A0(net232),
.A1(net240),
.A2(net237),
.A3(net233),
.S0(out17),
.S1(net649),
.X(net246)
);

sky130_fd_sc_hd__sdfsbp_2 c315(
.D(net231),
.SCD(net146),
.SCE(net121),
.SET_B(net142),
.CLK(clk),
.Q(net248),
.Q_N(net247)
);

sky130_fd_sc_hd__or4bb_4 c316(
.A(net237),
.B(net20),
.C_N(net245),
.D_N(net142),
.X(net249)
);

sky130_fd_sc_hd__a2111oi_4 c317(
.A1(net249),
.A2(net119),
.B1(out40),
.C1(net244),
.D1(net646),
.Y(net250)
);

sky130_fd_sc_hd__sdfxbp_1 c318(
.D(net150),
.SCD(net228),
.SCE(net250),
.CLK(clk),
.Q(net252),
.Q_N(net251)
);

sky130_fd_sc_hd__sdfxbp_2 c319(
.D(net250),
.SCD(out47),
.SCE(net252),
.CLK(clk),
.Q(net254),
.Q_N(net253)
);

sky130_fd_sc_hd__nor3_1 c320(
.A(net245),
.B(net248),
.C(out55),
.Y(net255)
);

sky130_fd_sc_hd__and3b_2 c321(
.A_N(net20),
.B(net84),
.C(net244),
.X(net256)
);

sky130_fd_sc_hd__sdfxtp_1 c322(
.D(net241),
.SCD(net215),
.SCE(net221),
.CLK(clk),
.Q(net257)
);

sky130_fd_sc_hd__nor3_1 c323(
.A(net255),
.B(net249),
.C(out55),
.Y(net258)
);

sky130_fd_sc_hd__sdfxtp_2 c324(
.D(net257),
.SCD(net146),
.SCE(net241),
.CLK(clk),
.Q(net259)
);

sky130_fd_sc_hd__or4bb_2 c325(
.A(net252),
.B(out1),
.C_N(net222),
.D_N(net142),
.X(net260)
);

sky130_fd_sc_hd__a2111oi_1 c326(
.A1(net259),
.A2(net260),
.B1(net253),
.C1(in17),
.D1(net142),
.Y(net261)
);

sky130_fd_sc_hd__sdfbbn_2 c327(
.D(net222),
.RESET_B(out40),
.SCD(net259),
.SCE(net261),
.SET_B(net257),
.CLK_N(clk),
.Q(out43),
.Q_N(net262)
);

sky130_fd_sc_hd__mux4_2 c328(
.A0(net258),
.A1(net228),
.A2(net257),
.A3(net260),
.S0(net145),
.S1(net220),
.X(net263)
);

sky130_fd_sc_hd__sdfbbp_1 c329(
.D(net260),
.RESET_B(net222),
.SCD(net18),
.SCE(net261),
.SET_B(out55),
.CLK(clk),
.Q(net265),
.Q_N(net264)
);

sky130_fd_sc_hd__mux4_2 c330(
.A0(net256),
.A1(net150),
.A2(net233),
.A3(net145),
.S0(net648),
.S1(net650),
.X(net266)
);

sky130_fd_sc_hd__sdfbbn_1 c331(
.D(net266),
.RESET_B(net8),
.SCD(net256),
.SCE(net264),
.SET_B(net261),
.CLK_N(clk),
.Q(net268),
.Q_N(net267)
);

sky130_fd_sc_hd__nand3_4 c332(
.A(net267),
.B(net260),
.C(net650),
.Y(net269)
);

sky130_fd_sc_hd__sdfbbn_2 c333(
.D(net268),
.RESET_B(net261),
.SCD(net254),
.SCE(net245),
.SET_B(net146),
.CLK_N(clk),
.Q(net271),
.Q_N(net270)
);

sky130_fd_sc_hd__mux4_4 c334(
.A0(net250),
.A1(net265),
.A2(net259),
.A3(net261),
.S0(net270),
.S1(net269),
.X(net272)
);

sky130_fd_sc_hd__mux4_2 c335(
.A0(net254),
.A1(net271),
.A2(net269),
.A3(net264),
.S0(in54),
.S1(out14),
.X(net273)
);

sky130_fd_sc_hd__and3_2 c336(
.A(net40),
.B(net271),
.C(out14),
.X(net274)
);

sky130_fd_sc_hd__sdfxtp_4 c337(
.D(net157),
.SCD(net164),
.SCE(net236),
.CLK(clk),
.Q(net275)
);

sky130_fd_sc_hd__nor3b_2 c338(
.A(net38),
.B(out51),
.C_N(net40),
.Y(net276)
);

sky130_fd_sc_hd__nand3_2 c339(
.A(net128),
.B(net275),
.C(net205),
.Y(out45)
);

sky130_fd_sc_hd__or3b_2 c340(
.A(net14),
.B(net274),
.C_N(in54),
.X(net277)
);

sky130_fd_sc_hd__nand3_1 c341(
.A(net146),
.B(net38),
.C(net251),
.Y(net278)
);

sky130_fd_sc_hd__mux4_1 c342(
.A0(net154),
.A1(net277),
.A2(net275),
.A3(net262),
.S0(out45),
.S1(net651),
.X(net279)
);

sky130_fd_sc_hd__nor3_4 c343(
.A(net277),
.B(net233),
.C(net275),
.Y(out61)
);

sky130_fd_sc_hd__dfbbn_1 c344(
.D(net164),
.RESET_B(net262),
.SET_B(out29),
.CLK_N(clk),
.Q(net281),
.Q_N(net280)
);

sky130_fd_sc_hd__sdfstp_1 c345(
.D(net121),
.SCD(net276),
.SCE(out40),
.SET_B(out17),
.CLK(clk),
.Q(net282)
);

sky130_fd_sc_hd__nand2b_1 c346(
.A_N(net274),
.B(net206),
.Y(out52)
);

sky130_fd_sc_hd__dfbbn_2 c347(
.D(net281),
.RESET_B(net275),
.SET_B(net238),
.CLK_N(clk),
.Q(net283)
);

sky130_fd_sc_hd__sdfstp_2 c348(
.D(net13),
.SCD(out61),
.SCE(net157),
.SET_B(out29),
.CLK(clk),
.Q(net284)
);

sky130_fd_sc_hd__dfbbp_1 c349(
.D(net246),
.RESET_B(out55),
.SET_B(net157),
.CLK(clk),
.Q(out32),
.Q_N(net285)
);

sky130_fd_sc_hd__and3b_2 c350(
.A_N(net145),
.B(net280),
.C(net282),
.X(net286)
);

sky130_fd_sc_hd__or4bb_1 c351(
.A(net159),
.B(net14),
.C_N(net284),
.D_N(net282),
.X(net287)
);

sky130_fd_sc_hd__or4bb_4 c352(
.A(net283),
.B(net284),
.C_N(net280),
.D_N(net119),
.X(net288)
);

sky130_fd_sc_hd__or4bb_2 c353(
.A(net155),
.B(net288),
.C_N(net159),
.D_N(net651),
.X(net289)
);

sky130_fd_sc_hd__mux4_2 c354(
.A0(net152),
.A1(net288),
.A2(net286),
.A3(net40),
.S0(net155),
.S1(net289),
.X(net290)
);

sky130_fd_sc_hd__sdfxbp_1 c355(
.D(net228),
.SCD(net290),
.SCE(net145),
.CLK(clk),
.Q(out27),
.Q_N(net291)
);

sky130_fd_sc_hd__mux4_4 c356(
.A0(net284),
.A1(in50),
.A2(net281),
.A3(out27),
.S0(net269),
.S1(net145),
.X(net292)
);

sky130_fd_sc_hd__mux4_2 c372(
.A0(net58),
.A1(net284),
.A2(out29),
.A3(out55),
.S0(in17),
.S1(out59),
.X(out48)
);

sky130_fd_sc_hd__mux4_4 c373(
.A0(in22),
.A1(net282),
.A2(net176),
.A3(out48),
.S0(out38),
.S1(net652),
.X(net293)
);

sky130_fd_sc_hd__mux4_2 c374(
.A0(net278),
.A1(net8),
.A2(out24),
.A3(out26),
.S0(out60),
.S1(net653),
.X(net294)
);

sky130_fd_sc_hd__mux4_2 c375(
.A0(in54),
.A1(out29),
.A2(net282),
.A3(out48),
.S0(net651),
.S1(out50),
.X(net295)
);

sky130_fd_sc_hd__mux4_1 c376(
.A0(net182),
.A1(out43),
.A2(net58),
.A3(out48),
.S0(net637),
.S1(out49),
.X(net296)
);

sky130_fd_sc_hd__mux4_1 c377(
.A0(net287),
.A1(net176),
.A2(net182),
.A3(out48),
.S0(out14),
.S1(out49),
.X(net297)
);

sky130_fd_sc_hd__nand2b_2 c378(
.A_N(net192),
.B(in14),
.Y(net298)
);

sky130_fd_sc_hd__nand2b_2 c379(
.A_N(net189),
.B(net200),
.Y(net299)
);

sky130_fd_sc_hd__dfrtn_1 c380(
.D(in9),
.RESET_B(net299),
.CLK_N(clk),
.Q(net300)
);

sky130_fd_sc_hd__dfrtp_1 c381(
.D(net299),
.RESET_B(net187),
.CLK(clk),
.Q(net301)
);

sky130_fd_sc_hd__and2_2 c382(
.A(net187),
.B(net184),
.X(net302)
);

sky130_fd_sc_hd__nand2b_1 c383(
.A_N(net195),
.B(net69),
.Y(net303)
);

sky130_fd_sc_hd__or3b_2 c384(
.A(net302),
.B(net301),
.C_N(net298),
.X(net304)
);

sky130_fd_sc_hd__and2b_1 c385(
.A_N(net185),
.B(net71),
.X(net305)
);

sky130_fd_sc_hd__nand3b_4 c386(
.A_N(net304),
.B(net298),
.C(net305),
.Y(net306)
);

sky130_fd_sc_hd__nor2_1 c387(
.A(net184),
.B(net305),
.Y(net307)
);

sky130_fd_sc_hd__or2b_1 c388(
.A(net305),
.B_N(net306),
.X(net308)
);

sky130_fd_sc_hd__nand2b_1 c389(
.A_N(net306),
.B(net71),
.Y(net309)
);

sky130_fd_sc_hd__nor3_4 c390(
.A(net194),
.B(net191),
.C(net303),
.Y(net310)
);

sky130_fd_sc_hd__or3_2 c391(
.A(net300),
.B(net305),
.C(out40),
.X(net311)
);

sky130_fd_sc_hd__a2111oi_1 c392(
.A1(net311),
.A2(net188),
.B1(net305),
.C1(net304),
.D1(net191),
.Y(net312)
);

sky130_fd_sc_hd__nor3b_1 c393(
.A(net312),
.B(net71),
.C_N(net305),
.Y(net313)
);

sky130_fd_sc_hd__sdfbbp_1 c394(
.D(net299),
.RESET_B(net300),
.SCD(net313),
.SCE(net71),
.SET_B(net308),
.CLK(clk),
.Q(net315),
.Q_N(net314)
);

sky130_fd_sc_hd__or3_2 c395(
.A(net200),
.B(net307),
.C(net313),
.X(net316)
);

sky130_fd_sc_hd__sdfstp_4 c396(
.D(net316),
.SCD(net313),
.SCE(net310),
.SET_B(net314),
.CLK(clk),
.Q(net317)
);

sky130_fd_sc_hd__sedfxbp_1 c397(
.D(net307),
.DE(net317),
.SCD(net298),
.SCE(net316),
.CLK(clk),
.Q(net319),
.Q_N(net318)
);

sky130_fd_sc_hd__nand2b_1 c398(
.A_N(net313),
.B(net201),
.Y(net320)
);

sky130_fd_sc_hd__or2b_2 c399(
.A(in30),
.B_N(net68),
.X(net321)
);

sky130_fd_sc_hd__or4bb_4 c400(
.A(in33),
.B(net212),
.C_N(net202),
.D_N(net221),
.X(net322)
);

sky130_fd_sc_hd__and2b_2 c401(
.A_N(net68),
.B(net302),
.X(net323)
);

sky130_fd_sc_hd__and2_1 c402(
.A(net311),
.B(net640),
.X(net324)
);

sky130_fd_sc_hd__or4bb_2 c403(
.A(net213),
.B(in36),
.C_N(net209),
.D_N(net640),
.X(net325)
);

sky130_fd_sc_hd__and3b_2 c404(
.A_N(net322),
.B(net307),
.C(net188),
.X(net326)
);

sky130_fd_sc_hd__mux4_2 c405(
.A0(in23),
.A1(net191),
.A2(net325),
.A3(net71),
.S0(net324),
.S1(net326),
.X(net327)
);

sky130_fd_sc_hd__nand3_2 c406(
.A(net323),
.B(net220),
.C(net326),
.Y(net328)
);

sky130_fd_sc_hd__a2111oi_4 c407(
.A1(net86),
.A2(net213),
.B1(net322),
.C1(net326),
.D1(out23),
.Y(net329)
);

sky130_fd_sc_hd__mux4_4 c408(
.A0(net328),
.A1(net68),
.A2(net221),
.A3(net326),
.S0(in30),
.S1(in27),
.X(net330)
);

sky130_fd_sc_hd__a2111oi_0 c409(
.A1(net306),
.A2(net327),
.B1(net324),
.C1(net326),
.D1(in17),
.Y(net331)
);

sky130_fd_sc_hd__sdfxbp_2 c410(
.D(net330),
.SCD(net326),
.SCE(net311),
.CLK(clk),
.Q(net333),
.Q_N(net332)
);

sky130_fd_sc_hd__sedfxbp_2 c411(
.D(net333),
.DE(net308),
.SCD(net331),
.SCE(net326),
.CLK(clk),
.Q(net335),
.Q_N(net334)
);

sky130_fd_sc_hd__or4bb_2 c412(
.A(net325),
.B(net220),
.C_N(net335),
.D_N(net326),
.X(net336)
);

sky130_fd_sc_hd__sdfxtp_1 c413(
.D(net331),
.SCD(net330),
.SCE(net326),
.CLK(clk),
.Q(net337)
);

sky130_fd_sc_hd__mux4_1 c414(
.A0(net335),
.A1(net298),
.A2(net221),
.A3(net84),
.S0(net326),
.S1(net332),
.X(net338)
);

sky130_fd_sc_hd__a2111o_2 c415(
.A1(net329),
.A2(net333),
.B1(net322),
.C1(net334),
.D1(net326),
.X(net339)
);

sky130_fd_sc_hd__sdfxtp_2 c416(
.D(net330),
.SCD(net337),
.SCE(net326),
.CLK(clk),
.Q(net340)
);

sky130_fd_sc_hd__sdfxtp_4 c417(
.D(net202),
.SCD(net339),
.SCE(net326),
.CLK(clk),
.Q(net341)
);

sky130_fd_sc_hd__sedfxtp_1 c418(
.D(net213),
.DE(net339),
.SCD(net325),
.SCE(net326),
.CLK(clk),
.Q(net342)
);

sky130_fd_sc_hd__or3_1 c419(
.A(net338),
.B(net342),
.C(net326),
.X(net343)
);

sky130_fd_sc_hd__nand3_2 c420(
.A(in39),
.B(net338),
.C(in33),
.Y(net344)
);

sky130_fd_sc_hd__sedfxtp_2 c421(
.D(net96),
.DE(net198),
.SCD(net339),
.SCE(net188),
.CLK(clk),
.Q(net345)
);

sky130_fd_sc_hd__and3_2 c422(
.A(net321),
.B(net236),
.C(net646),
.X(out30)
);

sky130_fd_sc_hd__sedfxtp_4 c423(
.D(net345),
.DE(net121),
.SCD(net191),
.SCE(net212),
.CLK(clk),
.Q(net346)
);

sky130_fd_sc_hd__or4bb_1 c424(
.A(net336),
.B(net206),
.C_N(in15),
.D_N(in54),
.X(net347)
);

sky130_fd_sc_hd__o2111ai_1 c425(
.A1(net341),
.A2(in39),
.B1(in54),
.C1(net234),
.D1(net326),
.Y(net348)
);

sky130_fd_sc_hd__or3b_1 c426(
.A(net327),
.B(net321),
.C_N(in54),
.X(net349)
);

sky130_fd_sc_hd__or3b_2 c427(
.A(net346),
.B(net336),
.C_N(net326),
.X(net350)
);

sky130_fd_sc_hd__mux4_2 c428(
.A0(net98),
.A1(net227),
.A2(net321),
.A3(net96),
.S0(net220),
.S1(net303),
.X(net351)
);

sky130_fd_sc_hd__sdfbbn_1 c429(
.D(net349),
.RESET_B(net212),
.SCD(net240),
.SCE(in61),
.SET_B(out17),
.CLK_N(clk),
.Q(net353),
.Q_N(net352)
);

sky130_fd_sc_hd__dfbbn_1 c430(
.D(net350),
.RESET_B(net128),
.SET_B(net323),
.CLK_N(clk),
.Q(net355),
.Q_N(net354)
);

sky130_fd_sc_hd__sdfrbp_1 c431(
.D(net348),
.RESET_B(net198),
.SCD(net350),
.SCE(net352),
.CLK(clk),
.Q(net357),
.Q_N(net356)
);

sky130_fd_sc_hd__sdfbbn_2 c432(
.D(net123),
.RESET_B(net234),
.SCD(net356),
.SCE(net238),
.SET_B(net355),
.CLK_N(clk),
.Q(net359),
.Q_N(net358)
);

sky130_fd_sc_hd__sdfbbp_1 c433(
.D(net357),
.RESET_B(in30),
.SCD(net347),
.SCE(net354),
.SET_B(net350),
.CLK(clk),
.Q(net361),
.Q_N(net360)
);

sky130_fd_sc_hd__or4bb_1 c434(
.A(net337),
.B(net355),
.C_N(net360),
.D_N(net96),
.X(net362)
);

sky130_fd_sc_hd__mux4_1 c435(
.A0(net298),
.A1(net357),
.A2(net353),
.A3(in39),
.S0(net119),
.S1(net112),
.X(out5)
);

sky130_fd_sc_hd__sdfrbp_2 c436(
.D(net344),
.RESET_B(net315),
.SCD(net355),
.SCE(out5),
.CLK(clk),
.Q(net364),
.Q_N(net363)
);

sky130_fd_sc_hd__a2111o_1 c437(
.A1(net355),
.A2(net364),
.B1(net352),
.C1(net188),
.D1(out5),
.X(net365)
);

sky130_fd_sc_hd__mux4_1 c438(
.A0(net364),
.A1(net346),
.A2(net356),
.A3(net354),
.S0(net365),
.S1(out5),
.X(net366)
);

sky130_fd_sc_hd__mux4_1 c439(
.A0(net227),
.A1(out5),
.A2(net366),
.A3(net317),
.S0(net356),
.S1(net354),
.X(net367)
);

sky130_fd_sc_hd__mux4_4 c440(
.A0(net347),
.A1(net366),
.A2(net357),
.A3(net351),
.S0(net310),
.S1(net363),
.X(net368)
);

sky130_fd_sc_hd__and2_1 c441(
.A(net353),
.B(net142),
.X(net369)
);

sky130_fd_sc_hd__or2b_1 c442(
.A(net359),
.B_N(in21),
.X(net370)
);

sky130_fd_sc_hd__nand3_2 c443(
.A(net255),
.B(net326),
.C(out5),
.Y(net371)
);

sky130_fd_sc_hd__sdfbbn_1 c444(
.D(net361),
.RESET_B(net364),
.SCD(net256),
.SCE(net358),
.SET_B(net339),
.CLK_N(clk),
.Q(net372)
);

sky130_fd_sc_hd__or2b_1 c445(
.A(net372),
.B_N(net370),
.X(net373)
);

sky130_fd_sc_hd__nand3b_4 c446(
.A_N(net369),
.B(net310),
.C(out5),
.Y(out37)
);

sky130_fd_sc_hd__nand3_1 c447(
.A(net373),
.B(net205),
.C(net370),
.Y(net374)
);

sky130_fd_sc_hd__o2111ai_2 c448(
.A1(net373),
.A2(net364),
.B1(net370),
.C1(net247),
.D1(out5),
.Y(net375)
);

sky130_fd_sc_hd__and3b_1 c449(
.A_N(net371),
.B(net365),
.C(net375),
.X(net376)
);

sky130_fd_sc_hd__nand2b_1 c450(
.A_N(net375),
.B(net363),
.Y(net377)
);

sky130_fd_sc_hd__or4bb_1 c451(
.A(net302),
.B(net255),
.C_N(net373),
.D_N(net370),
.X(net378)
);

sky130_fd_sc_hd__nand3_4 c452(
.A(net248),
.B(net370),
.C(net378),
.Y(net379)
);

sky130_fd_sc_hd__mux4_2 c453(
.A0(net378),
.A1(in56),
.A2(net373),
.A3(net375),
.S0(net142),
.S1(out5),
.X(net380)
);

sky130_fd_sc_hd__or3_1 c454(
.A(net377),
.B(net18),
.C(net378),
.X(net381)
);

sky130_fd_sc_hd__mux4_4 c455(
.A0(net376),
.A1(net261),
.A2(net18),
.A3(net375),
.S0(net378),
.S1(out17),
.X(net382)
);

sky130_fd_sc_hd__mux4_2 c456(
.A0(net374),
.A1(net378),
.A2(net363),
.A3(net379),
.S0(net381),
.S1(out17),
.X(net383)
);

sky130_fd_sc_hd__sdfbbn_2 c457(
.D(net261),
.RESET_B(net378),
.SCD(net142),
.SCE(net377),
.SET_B(net656),
.CLK_N(clk),
.Q(net385),
.Q_N(net384)
);

sky130_fd_sc_hd__mux4_2 c458(
.A0(net381),
.A1(net375),
.A2(net269),
.A3(net18),
.S0(net370),
.S1(net646),
.X(net386)
);

sky130_fd_sc_hd__mux4_1 c459(
.A0(in17),
.A1(net378),
.A2(net384),
.A3(net343),
.S0(net375),
.S1(net656),
.X(net387)
);

sky130_fd_sc_hd__o2111ai_1 c460(
.A1(net353),
.A2(net367),
.B1(out5),
.C1(net654),
.D1(net655),
.Y(net388)
);

sky130_fd_sc_hd__mux4_1 c461(
.A0(net388),
.A1(net339),
.A2(net378),
.A3(net238),
.S0(net384),
.S1(net655),
.X(net389)
);

sky130_fd_sc_hd__nor3b_2 c462(
.A(net362),
.B(out31),
.C_N(out45),
.Y(out15)
);

sky130_fd_sc_hd__mux4_1 c463(
.A0(net269),
.A1(net163),
.A2(net127),
.A3(out37),
.S0(in1),
.S1(out29),
.X(net390)
);

sky130_fd_sc_hd__mux4_2 c464(
.A0(net36),
.A1(out31),
.A2(net370),
.A3(out29),
.S0(net379),
.S1(net660),
.X(net391)
);

sky130_fd_sc_hd__mux4_1 c465(
.A0(net279),
.A1(net238),
.A2(out15),
.A3(net289),
.S0(in17),
.S1(net657),
.X(net392)
);

sky130_fd_sc_hd__sdfbbp_1 c466(
.D(net285),
.RESET_B(out15),
.SCD(net659),
.SCE(net661),
.SET_B(net663),
.CLK(clk),
.Q(net393)
);

sky130_fd_sc_hd__and3b_1 c467(
.A_N(net206),
.B(out42),
.C(net365),
.X(net394)
);

sky130_fd_sc_hd__and3b_4 c468(
.A_N(net271),
.B(net84),
.C(net663),
.X(net395)
);

sky130_fd_sc_hd__nand3b_1 c469(
.A_N(net270),
.B(net662),
.C(net663),
.Y(net396)
);

sky130_fd_sc_hd__mux4_1 c470(
.A0(net367),
.A1(out42),
.A2(net276),
.A3(net291),
.S0(net395),
.S1(out45),
.X(out9)
);

sky130_fd_sc_hd__mux4_2 c471(
.A0(net396),
.A1(net274),
.A2(net304),
.A3(net395),
.S0(net370),
.S1(net270),
.X(net397)
);

sky130_fd_sc_hd__and3_4 c472(
.A(net395),
.B(net304),
.C(net658),
.X(out46)
);

sky130_fd_sc_hd__and3_2 c473(
.A(net274),
.B(net291),
.C(net658),
.X(net398)
);

sky130_fd_sc_hd__and3b_1 c474(
.A_N(net317),
.B(net36),
.C(net310),
.X(out21)
);

sky130_fd_sc_hd__and3b_2 c475(
.A_N(net36),
.B(net303),
.C(net395),
.X(net399)
);

sky130_fd_sc_hd__mux4_4 c476(
.A0(net303),
.A1(net395),
.A2(net326),
.A3(net398),
.S0(out15),
.S1(out45),
.X(net400)
);

sky130_fd_sc_hd__nor3b_1 c477(
.A(net393),
.B(out21),
.C_N(out27),
.Y(net401)
);

sky130_fd_sc_hd__mux4_2 c478(
.A0(net399),
.A1(net365),
.A2(net34),
.A3(out9),
.S0(net84),
.S1(net661),
.X(net402)
);

sky130_fd_sc_hd__mux4_2 c479(
.A0(net401),
.A1(net286),
.A2(net395),
.A3(net279),
.S0(net398),
.S1(net663),
.X(net403)
);

sky130_fd_sc_hd__mux4_4 c480(
.A0(net397),
.A1(out5),
.A2(net395),
.A3(out9),
.S0(out15),
.S1(net665),
.X(net404)
);

sky130_fd_sc_hd__mux4_1 c481(
.A0(in50),
.A1(out37),
.A2(net395),
.A3(out15),
.S0(net667),
.S1(out41),
.X(net405)
);

sky130_fd_sc_hd__mux4_1 c482(
.A0(net395),
.A1(out29),
.A2(net36),
.A3(net34),
.S0(out41),
.S1(net668),
.X(net406)
);

sky130_fd_sc_hd__and2b_4 c504(
.A_N(net300),
.B(net318),
.X(net407)
);

sky130_fd_sc_hd__clkinv_2 c505(
.A(net636),
.Y(net408)
);

sky130_fd_sc_hd__nand2b_1 c506(
.A_N(in0),
.B(net408),
.Y(net409)
);

sky130_fd_sc_hd__nand2b_2 c507(
.A_N(net312),
.B(net69),
.Y(net410)
);

sky130_fd_sc_hd__dfbbn_2 c508(
.D(net316),
.RESET_B(net410),
.SET_B(net408),
.CLK_N(clk),
.Q(net412),
.Q_N(net411)
);

sky130_fd_sc_hd__nor2b_4 c509(
.A(net309),
.B_N(net412),
.Y(net413)
);

sky130_fd_sc_hd__buf_1 c510(
.A(net636),
.X(net414)
);

sky130_fd_sc_hd__a2111o_1 c511(
.A1(net407),
.A2(net408),
.B1(net413),
.C1(net414),
.D1(net410),
.X(net415)
);

sky130_fd_sc_hd__or2b_4 c512(
.A(net412),
.B_N(net408),
.X(net416)
);

sky130_fd_sc_hd__nand3b_2 c513(
.A_N(net201),
.B(net414),
.C(net188),
.Y(net417)
);

sky130_fd_sc_hd__and2b_4 c514(
.A_N(net410),
.B(net315),
.X(net418)
);

sky130_fd_sc_hd__nor3_4 c515(
.A(net416),
.B(net308),
.C(net415),
.Y(net419)
);

sky130_fd_sc_hd__dfrtp_2 c516(
.D(net419),
.RESET_B(net415),
.CLK(clk),
.Q(net420)
);

sky130_fd_sc_hd__nor3_2 c517(
.A(net409),
.B(net418),
.C(net414),
.Y(net421)
);

sky130_fd_sc_hd__nor2b_2 c518(
.A(net421),
.B_N(net414),
.Y(net422)
);

sky130_fd_sc_hd__dfbbp_1 c519(
.D(net407),
.RESET_B(net421),
.SET_B(net316),
.CLK(clk),
.Q(net424),
.Q_N(net423)
);

sky130_fd_sc_hd__sdfxbp_1 c520(
.D(net419),
.SCD(net422),
.SCE(net423),
.CLK(clk),
.Q(net426),
.Q_N(net425)
);

sky130_fd_sc_hd__mux4_2 c521(
.A0(net426),
.A1(net421),
.A2(net309),
.A3(net411),
.S0(net308),
.S1(net316),
.X(net427)
);

sky130_fd_sc_hd__sdfxbp_2 c522(
.D(net422),
.SCD(net424),
.SCE(net415),
.CLK(clk),
.Q(net429),
.Q_N(net428)
);

sky130_fd_sc_hd__mux4_4 c523(
.A0(net319),
.A1(net413),
.A2(net421),
.A3(net414),
.S0(net420),
.S1(net669),
.X(net430)
);

sky130_fd_sc_hd__mux4_1 c524(
.A0(net421),
.A1(net428),
.A2(net417),
.A3(net316),
.S0(net409),
.S1(net669),
.X(net431)
);

sky130_fd_sc_hd__nand3b_4 c525(
.A_N(net408),
.B(net188),
.C(net413),
.Y(net432)
);

sky130_fd_sc_hd__and3_1 c526(
.A(in14),
.B(net220),
.C(net432),
.X(net433)
);

sky130_fd_sc_hd__sdfxtp_1 c527(
.D(net414),
.SCD(net308),
.SCE(net430),
.CLK(clk),
.Q(net434)
);

sky130_fd_sc_hd__and3_4 c528(
.A(net429),
.B(net325),
.C(net434),
.X(net435)
);

sky130_fd_sc_hd__dfrtp_4 c529(
.D(in41),
.RESET_B(net430),
.CLK(clk),
.Q(net436)
);

sky130_fd_sc_hd__dfsbp_1 c530(
.D(net308),
.SET_B(net320),
.CLK(clk),
.Q(net438),
.Q_N(net437)
);

sky130_fd_sc_hd__and3b_1 c531(
.A_N(net432),
.B(net436),
.C(net670),
.X(net439)
);

sky130_fd_sc_hd__sdfxtp_2 c532(
.D(net71),
.SCD(net437),
.SCE(net343),
.CLK(clk),
.Q(net440)
);

sky130_fd_sc_hd__nor3b_1 c533(
.A(in17),
.B(net436),
.C_N(net71),
.Y(net441)
);

sky130_fd_sc_hd__sdfxtp_4 c534(
.D(net441),
.SCD(net439),
.SCE(net436),
.CLK(clk),
.Q(net442)
);

sky130_fd_sc_hd__dfbbn_1 c535(
.D(net436),
.RESET_B(net442),
.SET_B(net439),
.CLK_N(clk),
.Q(net444),
.Q_N(net443)
);

sky130_fd_sc_hd__dfbbn_2 c536(
.D(net430),
.RESET_B(net441),
.SET_B(net436),
.CLK_N(clk),
.Q(net445)
);

sky130_fd_sc_hd__or3b_2 c537(
.A(net435),
.B(net436),
.C_N(net85),
.X(net446)
);

sky130_fd_sc_hd__o2111a_1 c538(
.A1(net445),
.A2(net442),
.B1(net443),
.C1(net436),
.D1(net446),
.X(net447)
);

sky130_fd_sc_hd__o2111a_2 c539(
.A1(net324),
.A2(net85),
.B1(net440),
.C1(net446),
.D1(net188),
.X(net448)
);

sky130_fd_sc_hd__dfbbp_1 c540(
.D(net433),
.RESET_B(net446),
.SET_B(net444),
.CLK(clk),
.Q(net450),
.Q_N(net449)
);

sky130_fd_sc_hd__sdfbbn_1 c541(
.D(net305),
.RESET_B(net436),
.SCD(net448),
.SCE(net439),
.SET_B(net434),
.CLK_N(clk),
.Q(net452),
.Q_N(net451)
);

sky130_fd_sc_hd__a2111oi_1 c542(
.A1(net447),
.A2(net324),
.B1(net450),
.C1(net71),
.D1(net451),
.Y(out13)
);

sky130_fd_sc_hd__a2111o_2 c543(
.A1(net198),
.A2(net452),
.B1(net324),
.C1(out13),
.D1(net446),
.X(net453)
);

sky130_fd_sc_hd__sdfbbn_2 c544(
.D(net442),
.RESET_B(out13),
.SCD(net452),
.SCE(net450),
.SET_B(net453),
.CLK_N(clk),
.Q(net454)
);

sky130_fd_sc_hd__sdfbbp_1 c545(
.D(net454),
.RESET_B(net453),
.SCD(net339),
.SCE(net438),
.SET_B(net451),
.CLK(clk),
.Q(net456),
.Q_N(net455)
);

sky130_fd_sc_hd__sdfxbp_1 c546(
.D(net438),
.SCD(net343),
.SCE(net112),
.CLK(clk),
.Q(net458),
.Q_N(net457)
);

sky130_fd_sc_hd__and3b_1 c547(
.A_N(in50),
.B(in27),
.C(net365),
.X(net459)
);

sky130_fd_sc_hd__sdfbbn_1 c548(
.D(net458),
.RESET_B(net85),
.SCD(net417),
.SCE(net459),
.SET_B(net440),
.CLK_N(clk),
.Q(net461),
.Q_N(net460)
);

sky130_fd_sc_hd__or3_1 c549(
.A(net461),
.B(net452),
.C(net434),
.X(net462)
);

sky130_fd_sc_hd__mux4_2 c550(
.A0(net240),
.A1(net462),
.A2(net434),
.A3(net451),
.S0(out13),
.S1(net112),
.X(net463)
);

sky130_fd_sc_hd__mux4_1 c551(
.A0(net440),
.A1(net351),
.A2(net338),
.A3(net449),
.S0(net459),
.S1(net339),
.X(net464)
);

sky130_fd_sc_hd__a2111oi_4 c552(
.A1(net234),
.A2(out13),
.B1(net459),
.C1(net437),
.D1(net460),
.Y(net465)
);

sky130_fd_sc_hd__sdfbbn_2 c553(
.D(net465),
.RESET_B(net412),
.SCD(net461),
.SCE(net314),
.SET_B(net671),
.CLK_N(clk),
.Q(net467),
.Q_N(net466)
);

sky130_fd_sc_hd__sdfbbp_1 c554(
.D(net221),
.RESET_B(net112),
.SCD(net351),
.SCE(net465),
.SET_B(net671),
.CLK(clk),
.Q(net468)
);

sky130_fd_sc_hd__sdfbbn_1 c555(
.D(in27),
.RESET_B(net112),
.SCD(net466),
.SCE(net465),
.SET_B(net671),
.CLK_N(clk),
.Q(net470),
.Q_N(net469)
);

sky130_fd_sc_hd__sdfxbp_2 c556(
.D(net467),
.SCD(net417),
.SCE(net342),
.CLK(clk),
.Q(out19),
.Q_N(net471)
);

sky130_fd_sc_hd__o2111a_2 c557(
.A1(net459),
.A2(net434),
.B1(out19),
.C1(net469),
.D1(out5),
.X(net472)
);

sky130_fd_sc_hd__mux4_1 c558(
.A0(net470),
.A1(net365),
.A2(net465),
.A3(net412),
.S0(net463),
.S1(net471),
.X(net473)
);

sky130_fd_sc_hd__mux4_4 c559(
.A0(net472),
.A1(net85),
.A2(in0),
.A3(net669),
.S0(net671),
.S1(net672),
.X(net474)
);

sky130_fd_sc_hd__mux4_2 c560(
.A0(net188),
.A1(net474),
.A2(net465),
.A3(net457),
.S0(net669),
.S1(net672),
.X(net475)
);

sky130_fd_sc_hd__a2111oi_2 c561(
.A1(net468),
.A2(out19),
.B1(net450),
.C1(net474),
.D1(net672),
.Y(net476)
);

sky130_fd_sc_hd__mux4_4 c562(
.A0(net474),
.A1(net338),
.A2(net459),
.A3(net471),
.S0(net476),
.S1(net672),
.X(net477)
);

sky130_fd_sc_hd__mux4_4 c563(
.A0(net476),
.A1(net459),
.A2(net474),
.A3(net351),
.S0(net471),
.S1(net675),
.X(net478)
);

sky130_fd_sc_hd__mux4_4 c564(
.A0(net315),
.A1(net338),
.A2(net411),
.A3(net474),
.S0(net673),
.S1(net674),
.X(net479)
);

sky130_fd_sc_hd__mux4_1 c565(
.A0(net479),
.A1(net472),
.A2(out19),
.A3(net474),
.S0(net465),
.S1(net675),
.X(net480)
);

sky130_fd_sc_hd__mux4_1 c566(
.A0(out1),
.A1(net479),
.A2(in56),
.A3(net674),
.S0(net677),
.S1(net678),
.X(net481)
);

sky130_fd_sc_hd__sdfbbn_2 c567(
.D(net351),
.RESET_B(net444),
.SCD(net265),
.SCE(net420),
.SET_B(net339),
.CLK_N(clk),
.Q(net483),
.Q_N(net482)
);

sky130_fd_sc_hd__or3b_1 c568(
.A(net18),
.B(out19),
.C_N(out17),
.X(net484)
);

sky130_fd_sc_hd__mux4_1 c569(
.A0(net484),
.A1(net385),
.A2(out1),
.A3(net18),
.S0(net443),
.S1(out13),
.X(net485)
);

sky130_fd_sc_hd__sdfbbp_1 c570(
.D(net265),
.RESET_B(net343),
.SCD(net142),
.SCE(net339),
.SET_B(out5),
.CLK(clk),
.Q(net487),
.Q_N(net486)
);

sky130_fd_sc_hd__mux4_4 c571(
.A0(net339),
.A1(net448),
.A2(net119),
.A3(net142),
.S0(net379),
.S1(net482),
.X(net488)
);

sky130_fd_sc_hd__mux4_2 c572(
.A0(net484),
.A1(net142),
.A2(net370),
.A3(net448),
.S0(net676),
.S1(net680),
.X(net489)
);

sky130_fd_sc_hd__nor3b_1 c573(
.A(net265),
.B(net677),
.C_N(net680),
.Y(net490)
);

sky130_fd_sc_hd__mux4_4 c574(
.A0(net487),
.A1(net256),
.A2(net455),
.A3(net489),
.S0(net85),
.S1(out5),
.X(net491)
);

sky130_fd_sc_hd__a2111o_1 c575(
.A1(net342),
.A2(net486),
.B1(net490),
.C1(out5),
.D1(net448),
.X(net492)
);

sky130_fd_sc_hd__or4bb_4 c576(
.A(net490),
.B(net342),
.C_N(net492),
.D_N(out5),
.X(net493)
);

sky130_fd_sc_hd__sdfxtp_1 c577(
.D(net485),
.SCD(net351),
.SCE(net448),
.CLK(clk),
.Q(net494)
);

sky130_fd_sc_hd__mux4_4 c578(
.A0(net212),
.A1(net343),
.A2(net494),
.A3(net482),
.S0(net455),
.S1(net476),
.X(net495)
);

sky130_fd_sc_hd__or4bb_4 c579(
.A(net494),
.B(net448),
.C_N(in17),
.D_N(net326),
.X(net496)
);

sky130_fd_sc_hd__mux4_4 c580(
.A0(net493),
.A1(net492),
.A2(net264),
.A3(net384),
.S0(net142),
.S1(net679),
.X(net497)
);

sky130_fd_sc_hd__or3_1 c581(
.A(net492),
.B(net310),
.C(net342),
.X(net498)
);

sky130_fd_sc_hd__mux4_4 c582(
.A0(net491),
.A1(out13),
.A2(net492),
.A3(net351),
.S0(net483),
.S1(net493),
.X(net499)
);

sky130_fd_sc_hd__mux4_1 c583(
.A0(net380),
.A1(in15),
.A2(net491),
.A3(net496),
.S0(net448),
.S1(net142),
.X(net500)
);

sky130_fd_sc_hd__mux4_4 c584(
.A0(net448),
.A1(net142),
.A2(net471),
.A3(net84),
.S0(net683),
.S1(net686),
.X(net501)
);

sky130_fd_sc_hd__mux4_2 c585(
.A0(net498),
.A1(net501),
.A2(net420),
.A3(net379),
.S0(net492),
.S1(net683),
.X(net502)
);

sky130_fd_sc_hd__mux4_1 c586(
.A0(net501),
.A1(net142),
.A2(out17),
.A3(out14),
.S0(net680),
.S1(net685),
.X(net503)
);

sky130_fd_sc_hd__mux4_2 c587(
.A0(net264),
.A1(out14),
.A2(net679),
.A3(net680),
.S0(net681),
.S1(net687),
.X(net504)
);

sky130_fd_sc_hd__mux4_4 c588(
.A0(net420),
.A1(net385),
.A2(net490),
.A3(net288),
.S0(out5),
.S1(net684),
.X(net505)
);

sky130_fd_sc_hd__mux4_1 c589(
.A0(net505),
.A1(net398),
.A2(net289),
.A3(net385),
.S0(net34),
.S1(net394),
.X(net506)
);

sky130_fd_sc_hd__mux4_2 c590(
.A0(net394),
.A1(net34),
.A2(net365),
.A3(net504),
.S0(out15),
.S1(net482),
.X(net507)
);

sky130_fd_sc_hd__mux4_1 c591(
.A0(net448),
.A1(net412),
.A2(net163),
.A3(net34),
.S0(net504),
.S1(net326),
.X(net508)
);

sky130_fd_sc_hd__mux4_2 c592(
.A0(net490),
.A1(net379),
.A2(net326),
.A3(out15),
.S0(net679),
.S1(net688),
.X(net509)
);

sky130_fd_sc_hd__mux4_2 c593(
.A0(net462),
.A1(net506),
.A2(net394),
.A3(net163),
.S0(net288),
.S1(net476),
.X(net510)
);

sky130_fd_sc_hd__mux4_2 c594(
.A0(in61),
.A1(net310),
.A2(net412),
.A3(net34),
.S0(out21),
.S1(net681),
.X(net511)
);

sky130_fd_sc_hd__mux4_2 c595(
.A0(net84),
.A1(net504),
.A2(in17),
.A3(net664),
.S0(net687),
.S1(net688),
.X(net512)
);

sky130_fd_sc_hd__mux4_1 c596(
.A0(net85),
.A1(out1),
.A2(net289),
.A3(net304),
.S0(net688),
.S1(net689),
.X(net513)
);

sky130_fd_sc_hd__mux4_1 c597(
.A0(net406),
.A1(net370),
.A2(net398),
.A3(net304),
.S0(net664),
.S1(net666),
.X(net514)
);

sky130_fd_sc_hd__mux4_4 c598(
.A0(net512),
.A1(net84),
.A2(net514),
.A3(net289),
.S0(out14),
.S1(net684),
.X(net515)
);

sky130_fd_sc_hd__mux4_1 c599(
.A0(net514),
.A1(net398),
.A2(net34),
.A3(net163),
.S0(net370),
.S1(net411),
.X(net516)
);

sky130_fd_sc_hd__mux4_4 c600(
.A0(net365),
.A1(net288),
.A2(net289),
.A3(net511),
.S0(net482),
.S1(net690),
.X(net517)
);

sky130_fd_sc_hd__mux4_2 c601(
.A0(net163),
.A1(net288),
.A2(net398),
.A3(out13),
.S0(net84),
.S1(net688),
.X(out25)
);

sky130_fd_sc_hd__mux4_2 c602(
.A0(net310),
.A1(net511),
.A2(net163),
.A3(out15),
.S0(net365),
.S1(net681),
.X(net518)
);

sky130_fd_sc_hd__mux4_2 c603(
.A0(out15),
.A1(net411),
.A2(out17),
.A3(net690),
.S0(net691),
.S1(net693),
.X(net519)
);

sky130_fd_sc_hd__mux4_1 c604(
.A0(net220),
.A1(in61),
.A2(net513),
.A3(net684),
.S0(net689),
.S1(net694),
.X(net520)
);

sky130_fd_sc_hd__mux4_1 c605(
.A0(net517),
.A1(net504),
.A2(net514),
.A3(out1),
.S0(net694),
.S1(net695),
.X(net521)
);

sky130_fd_sc_hd__mux4_1 c606(
.A0(net452),
.A1(net119),
.A2(out14),
.A3(net687),
.S0(net688),
.S1(net692),
.X(net522)
);

sky130_fd_sc_hd__mux4_2 c607(
.A0(net119),
.A1(out9),
.A2(net513),
.A3(net511),
.S0(in17),
.S1(net696),
.X(net523)
);

sky130_fd_sc_hd__mux4_4 c608(
.A0(net522),
.A1(net411),
.A2(net688),
.A3(net689),
.S0(out11),
.S1(net698),
.X(out22)
);

sky130_fd_sc_hd__or2_1 c630(
.A(net69),
.B(net409),
.X(net524)
);

sky130_fd_sc_hd__and2_4 c631(
.A(net416),
.B(net69),
.X(net525)
);

sky130_fd_sc_hd__and3b_1 c632(
.A_N(net186),
.B(net409),
.C(net524),
.X(net526)
);

sky130_fd_sc_hd__and2b_4 c633(
.A_N(net424),
.B(net410),
.X(out4)
);

sky130_fd_sc_hd__nor3b_2 c634(
.A(net526),
.B(net409),
.C_N(out4),
.Y(net527)
);

sky130_fd_sc_hd__or4bb_2 c635(
.A(net410),
.B(net525),
.C_N(net186),
.D_N(out4),
.X(net528)
);

sky130_fd_sc_hd__and3_2 c636(
.A(net525),
.B(net425),
.C(out4),
.X(net529)
);

sky130_fd_sc_hd__or4bb_1 c637(
.A(net529),
.B(net528),
.C_N(net413),
.D_N(net670),
.X(net530)
);

sky130_fd_sc_hd__and3_2 c638(
.A(net524),
.B(net186),
.C(net525),
.X(net531)
);

sky130_fd_sc_hd__or4bb_2 c639(
.A(net531),
.B(net525),
.C_N(net527),
.D_N(net409),
.X(net532)
);

sky130_fd_sc_hd__nor3_1 c640(
.A(net528),
.B(net301),
.C(in17),
.Y(net533)
);

sky130_fd_sc_hd__dfsbp_2 c641(
.D(net532),
.SET_B(net528),
.CLK(clk),
.Q(net535),
.Q_N(net534)
);

sky130_fd_sc_hd__sdfxtp_2 c642(
.D(net415),
.SCD(net531),
.SCE(net530),
.CLK(clk),
.Q(net536)
);

sky130_fd_sc_hd__nor2b_1 c643(
.A(net426),
.B_N(net527),
.Y(net537)
);

sky130_fd_sc_hd__sdfrtn_1 c644(
.D(net533),
.RESET_B(net535),
.SCD(net527),
.SCE(net69),
.CLK_N(clk),
.Q(net538)
);

sky130_fd_sc_hd__sdfxtp_4 c645(
.D(net418),
.SCD(net530),
.SCE(out4),
.CLK(clk),
.Q(net539)
);

sky130_fd_sc_hd__dfbbn_1 c646(
.D(net537),
.RESET_B(net533),
.SET_B(net526),
.CLK_N(clk),
.Q(net541),
.Q_N(net540)
);

sky130_fd_sc_hd__sdfrtp_1 c647(
.D(net532),
.RESET_B(net538),
.SCD(net536),
.SCE(net524),
.CLK(clk),
.Q(net542)
);

sky130_fd_sc_hd__mux4_2 c648(
.A0(net542),
.A1(net527),
.A2(net540),
.A3(net410),
.S0(net534),
.S1(net524),
.X(net543)
);

sky130_fd_sc_hd__mux4_1 c649(
.A0(net541),
.A1(net536),
.A2(net537),
.A3(net301),
.S0(net543),
.S1(net539),
.X(net544)
);

sky130_fd_sc_hd__mux4_2 c650(
.A0(net538),
.A1(net524),
.A2(net542),
.A3(net543),
.S0(net410),
.S1(net531),
.X(net545)
);

sky130_fd_sc_hd__sdfrtp_2 c651(
.D(net209),
.RESET_B(net528),
.SCD(net417),
.SCE(net420),
.CLK(clk),
.Q(net546)
);

sky130_fd_sc_hd__or3b_2 c652(
.A(net340),
.B(net449),
.C_N(net670),
.X(net547)
);

sky130_fd_sc_hd__nand2b_2 c653(
.A_N(net340),
.B(net536),
.Y(net548)
);

sky130_fd_sc_hd__dfbbn_2 c654(
.D(net320),
.RESET_B(net221),
.SET_B(net699),
.CLK_N(clk),
.Q(net550),
.Q_N(net549)
);

sky130_fd_sc_hd__dfbbp_1 c655(
.D(net413),
.RESET_B(net526),
.SET_B(net543),
.CLK(clk),
.Q(net551)
);

sky130_fd_sc_hd__sdfrtp_4 c656(
.D(net530),
.RESET_B(net320),
.SCD(net546),
.SCE(net550),
.CLK(clk),
.Q(net552)
);

sky130_fd_sc_hd__nand3b_1 c657(
.A_N(net546),
.B(net456),
.C(net534),
.Y(net553)
);

sky130_fd_sc_hd__or4bb_1 c658(
.A(in16),
.B(net221),
.C_N(net528),
.D_N(net699),
.X(net554)
);

sky130_fd_sc_hd__mux4_4 c659(
.A0(net553),
.A1(net552),
.A2(net546),
.A3(net340),
.S0(net529),
.S1(net699),
.X(net555)
);

sky130_fd_sc_hd__mux4_2 c660(
.A0(net550),
.A1(net543),
.A2(net547),
.A3(out23),
.S0(out3),
.S1(net699),
.X(net556)
);

sky130_fd_sc_hd__nor3b_4 c661(
.A(in16),
.B(net548),
.C_N(net209),
.Y(net557)
);

sky130_fd_sc_hd__nor3b_2 c662(
.A(net301),
.B(net420),
.C_N(net413),
.Y(net558)
);

sky130_fd_sc_hd__sdfxbp_1 c663(
.D(net543),
.SCD(net301),
.SCE(net554),
.CLK(clk),
.Q(net559)
);

sky130_fd_sc_hd__sdfsbp_1 c664(
.D(net453),
.SCD(net557),
.SCE(out4),
.SET_B(net700),
.CLK(clk),
.Q(net561),
.Q_N(net560)
);

sky130_fd_sc_hd__a2111oi_2 c665(
.A1(net529),
.A2(net552),
.B1(net549),
.C1(net557),
.D1(net700),
.Y(net562)
);

sky130_fd_sc_hd__sdfsbp_2 c666(
.D(net551),
.SCD(net530),
.SCE(net449),
.SET_B(net699),
.CLK(clk),
.Q(net563)
);

sky130_fd_sc_hd__sdfstp_1 c667(
.D(net559),
.SCD(net320),
.SCE(net554),
.SET_B(net340),
.CLK(clk),
.Q(net564)
);

sky130_fd_sc_hd__or3b_2 c668(
.A(net561),
.B(net564),
.C_N(net548),
.X(net565)
);

sky130_fd_sc_hd__sdfstp_2 c669(
.D(net562),
.SCD(net564),
.SCE(net546),
.SET_B(net670),
.CLK(clk),
.Q(net566)
);

sky130_fd_sc_hd__nor3_2 c670(
.A(net558),
.B(net565),
.C(net564),
.Y(net567)
);

sky130_fd_sc_hd__or4bb_4 c671(
.A(net563),
.B(net548),
.C_N(net546),
.D_N(out3),
.X(net568)
);

sky130_fd_sc_hd__sdfbbn_1 c672(
.D(net112),
.RESET_B(net420),
.SCD(net463),
.SCE(net530),
.SET_B(net669),
.CLK_N(clk),
.Q(net570),
.Q_N(net569)
);

sky130_fd_sc_hd__mux4_2 c673(
.A0(net555),
.A1(out4),
.A2(net450),
.A3(net539),
.S0(net420),
.S1(net671),
.X(net571)
);

sky130_fd_sc_hd__sdfbbn_2 c674(
.D(net552),
.RESET_B(net539),
.SCD(net476),
.SCE(net569),
.SET_B(net669),
.CLK_N(clk),
.Q(net573),
.Q_N(net572)
);

sky130_fd_sc_hd__mux4_4 c675(
.A0(net570),
.A1(net539),
.A2(net420),
.A3(net567),
.S0(net547),
.S1(out3),
.X(net574)
);

sky130_fd_sc_hd__sdfbbp_1 c676(
.D(net573),
.RESET_B(in33),
.SCD(net476),
.SCE(net455),
.SET_B(net672),
.CLK(clk),
.Q(net576),
.Q_N(net575)
);

sky130_fd_sc_hd__a2111oi_1 c677(
.A1(net525),
.A2(net561),
.B1(net547),
.C1(net539),
.D1(out5),
.Y(net577)
);

sky130_fd_sc_hd__mux4_1 c678(
.A0(net557),
.A1(net569),
.A2(net112),
.A3(net575),
.S0(net672),
.S1(net702),
.X(net578)
);

sky130_fd_sc_hd__mux4_4 c679(
.A0(net463),
.A1(net450),
.A2(net570),
.A3(net560),
.S0(net525),
.S1(in5),
.X(net579)
);

sky130_fd_sc_hd__a2111o_2 c680(
.A1(net552),
.A2(net576),
.B1(net547),
.C1(net577),
.D1(net112),
.X(out0)
);

sky130_fd_sc_hd__a2111o_4 c681(
.A1(net576),
.A2(net85),
.B1(out5),
.C1(net671),
.D1(net672),
.X(net580)
);

sky130_fd_sc_hd__sdfbbn_1 c682(
.D(net539),
.RESET_B(net554),
.SCD(net573),
.SCE(net566),
.SET_B(net646),
.CLK_N(clk),
.Q(net581)
);

sky130_fd_sc_hd__sdfbbn_2 c683(
.D(net417),
.RESET_B(net238),
.SCD(out4),
.SCE(net463),
.SET_B(net569),
.CLK_N(clk),
.Q(net583),
.Q_N(net582)
);

sky130_fd_sc_hd__mux4_2 c684(
.A0(net191),
.A1(net567),
.A2(net582),
.A3(out4),
.S0(net547),
.S1(net417),
.X(net584)
);

sky130_fd_sc_hd__mux4_1 c685(
.A0(net577),
.A1(net580),
.A2(net570),
.A3(net582),
.S0(net220),
.S1(net575),
.X(net585)
);

sky130_fd_sc_hd__a2111o_2 c686(
.A1(net583),
.A2(net561),
.B1(net585),
.C1(net573),
.D1(net575),
.X(net586)
);

sky130_fd_sc_hd__a2111oi_2 c687(
.A1(net581),
.A2(in56),
.B1(net576),
.C1(in33),
.D1(net704),
.Y(net587)
);

sky130_fd_sc_hd__mux4_4 c688(
.A0(net587),
.A1(net578),
.A2(net567),
.A3(net417),
.S0(net449),
.S1(net672),
.X(net588)
);

sky130_fd_sc_hd__mux4_2 c689(
.A0(net547),
.A1(out5),
.A2(net566),
.A3(out0),
.S0(net560),
.S1(net701),
.X(net589)
);

sky130_fd_sc_hd__sdfbbp_1 c690(
.D(net583),
.RESET_B(out4),
.SCD(net417),
.SCE(net703),
.SET_B(net705),
.CLK(clk),
.Q(net590)
);

sky130_fd_sc_hd__mux4_2 c691(
.A0(net589),
.A1(net590),
.A2(net238),
.A3(net572),
.S0(in56),
.S1(net669),
.X(net591)
);

sky130_fd_sc_hd__o2111a_4 c692(
.A1(net527),
.A2(net191),
.B1(net314),
.C1(net705),
.D1(net706),
.X(net592)
);

sky130_fd_sc_hd__a2111oi_4 c693(
.A1(net564),
.A2(net536),
.B1(in36),
.C1(in56),
.D1(in17),
.Y(net593)
);

sky130_fd_sc_hd__sdfbbn_1 c694(
.D(net578),
.RESET_B(net592),
.SCD(net483),
.SCE(net585),
.SET_B(net326),
.CLK_N(clk),
.Q(net595),
.Q_N(net594)
);

sky130_fd_sc_hd__mux4_4 c695(
.A0(net585),
.A1(out5),
.A2(net535),
.A3(net594),
.S0(net142),
.S1(net326),
.X(net596)
);

sky130_fd_sc_hd__mux4_4 c696(
.A0(net304),
.A1(net586),
.A2(net595),
.A3(net585),
.S0(net256),
.S1(net682),
.X(net597)
);

sky130_fd_sc_hd__mux4_2 c697(
.A0(net256),
.A1(in36),
.A2(net476),
.A3(out5),
.S0(out14),
.S1(net703),
.X(net598)
);

sky130_fd_sc_hd__mux4_2 c698(
.A0(net343),
.A1(net593),
.A2(in11),
.A3(in17),
.S0(net703),
.S1(net704),
.X(net599)
);

sky130_fd_sc_hd__mux4_2 c699(
.A0(net595),
.A1(net85),
.A2(out5),
.A3(in17),
.S0(out14),
.S1(net704),
.X(net600)
);

sky130_fd_sc_hd__mux4_1 c700(
.A0(net597),
.A1(in21),
.A2(net586),
.A3(net379),
.S0(net343),
.S1(net703),
.X(net601)
);

sky130_fd_sc_hd__o2111a_4 c701(
.A1(net315),
.A2(net600),
.B1(net566),
.C1(net142),
.D1(net568),
.X(net602)
);

sky130_fd_sc_hd__mux4_2 c702(
.A0(net535),
.A1(out0),
.A2(net476),
.A3(net564),
.S0(net142),
.S1(net671),
.X(net603)
);

sky130_fd_sc_hd__sdfbbn_2 c703(
.D(net142),
.RESET_B(net476),
.SCD(net420),
.SCE(net671),
.SET_B(net708),
.CLK_N(clk),
.Q(out2),
.Q_N(net604)
);

sky130_fd_sc_hd__mux4_1 c704(
.A0(net536),
.A1(net503),
.A2(net220),
.A3(net384),
.S0(net476),
.S1(net526),
.X(net605)
);

sky130_fd_sc_hd__mux4_1 c705(
.A0(net385),
.A1(net256),
.A2(in17),
.A3(net572),
.S0(net712),
.S1(net714),
.X(net606)
);

sky130_fd_sc_hd__a2111oi_2 c706(
.A1(net606),
.A2(net142),
.B1(net708),
.C1(net709),
.D1(net711),
.Y(net607)
);

sky130_fd_sc_hd__mux4_2 c707(
.A0(net573),
.A1(net503),
.A2(net600),
.A3(in17),
.S0(net455),
.S1(net710),
.X(net608)
);

sky130_fd_sc_hd__sdfbbp_1 c708(
.D(net596),
.RESET_B(net592),
.SCD(out5),
.SCE(net704),
.SET_B(net713),
.CLK(clk),
.Q(net609)
);

sky130_fd_sc_hd__a2111o_1 c709(
.A1(net593),
.A2(net607),
.B1(net326),
.C1(out0),
.D1(net596),
.X(net610)
);

sky130_fd_sc_hd__mux4_2 c710(
.A0(net602),
.A1(net593),
.A2(out1),
.A3(net238),
.S0(net572),
.S1(net682),
.X(net611)
);

sky130_fd_sc_hd__mux4_4 c711(
.A0(net526),
.A1(net600),
.A2(net142),
.A3(net566),
.S0(net597),
.S1(net710),
.X(net612)
);

sky130_fd_sc_hd__mux4_4 c712(
.A0(net566),
.A1(net610),
.A2(in56),
.A3(net220),
.S0(net700),
.S1(net715),
.X(net613)
);

sky130_fd_sc_hd__sdfbbn_1 c713(
.D(out0),
.RESET_B(net610),
.SCD(net712),
.SCE(net714),
.SET_B(net718),
.CLK_N(clk),
.Q(net614)
);

sky130_fd_sc_hd__mux4_1 c714(
.A0(net34),
.A1(net289),
.A2(out1),
.A3(net456),
.S0(in0),
.S1(net707),
.X(net615)
);

sky130_fd_sc_hd__mux4_2 c715(
.A0(net238),
.A1(net615),
.A2(net483),
.A3(in21),
.S0(net455),
.S1(net698),
.X(net616)
);

sky130_fd_sc_hd__mux4_1 c716(
.A0(net508),
.A1(net398),
.A2(net238),
.A3(net615),
.S0(out3),
.S1(net719),
.X(net617)
);

sky130_fd_sc_hd__mux4_1 c717(
.A0(net456),
.A1(net496),
.A2(in17),
.A3(out4),
.S0(out1),
.S1(net716),
.X(net618)
);

sky130_fd_sc_hd__mux4_2 c718(
.A0(net609),
.A1(net276),
.A2(net496),
.A3(out23),
.S0(net691),
.S1(net700),
.X(net619)
);

sky130_fd_sc_hd__mux4_1 c719(
.A0(net221),
.A1(net85),
.A2(net604),
.A3(net511),
.S0(net698),
.S1(net720),
.X(net620)
);

sky130_fd_sc_hd__mux4_2 c720(
.A0(net511),
.A1(net615),
.A2(net619),
.A3(out5),
.S0(out1),
.S1(out14),
.X(net621)
);

sky130_fd_sc_hd__mux4_1 c721(
.A0(net496),
.A1(net398),
.A2(out0),
.A3(net697),
.S0(net700),
.S1(net719),
.X(net622)
);

sky130_fd_sc_hd__mux4_4 c722(
.A0(net614),
.A1(net610),
.A2(out5),
.A3(net379),
.S0(out4),
.S1(net420),
.X(net623)
);

sky130_fd_sc_hd__mux4_2 c723(
.A0(net513),
.A1(net489),
.A2(out0),
.A3(net34),
.S0(net691),
.S1(net707),
.X(net624)
);

sky130_fd_sc_hd__mux4_2 c724(
.A0(net483),
.A1(net513),
.A2(net489),
.A3(net326),
.S0(out0),
.S1(net691),
.X(net625)
);

sky130_fd_sc_hd__mux4_2 c725(
.A0(net568),
.A1(net622),
.A2(net379),
.A3(net385),
.S0(net420),
.S1(net456),
.X(net626)
);

sky130_fd_sc_hd__mux4_1 c726(
.A0(net276),
.A1(net476),
.A2(net85),
.A3(net34),
.S0(net722),
.S1(net723),
.X(net627)
);

sky130_fd_sc_hd__mux4_2 c727(
.A0(net326),
.A1(out0),
.A2(in56),
.A3(net698),
.S0(net717),
.S1(net721),
.X(net628)
);

sky130_fd_sc_hd__mux4_1 c728(
.A0(net620),
.A1(out0),
.A2(out1),
.A3(net398),
.S0(net723),
.S1(net724),
.X(net629)
);

sky130_fd_sc_hd__mux4_2 c729(
.A0(net379),
.A1(net619),
.A2(net398),
.A3(net289),
.S0(net238),
.S1(net725),
.X(net630)
);

sky130_fd_sc_hd__mux4_2 c730(
.A0(in21),
.A1(net511),
.A2(net707),
.A3(net726),
.S0(net727),
.S1(net728),
.X(net631)
);

sky130_fd_sc_hd__mux4_1 c731(
.A0(net476),
.A1(net631),
.A2(in56),
.A3(net722),
.S0(net723),
.S1(net726),
.X(net632)
);

sky130_fd_sc_hd__mux4_2 c732(
.A0(net631),
.A1(out0),
.A2(net238),
.A3(net719),
.S0(net726),
.S1(net729),
.X(net633)
);

sky130_fd_sc_hd__mux4_1 c733(
.A0(net370),
.A1(net618),
.A2(net628),
.A3(out0),
.S0(out1),
.S1(net631),
.X(net634)
);

sky130_fd_sc_hd__mux4_4 c734(
.A0(net489),
.A1(net456),
.A2(net631),
.A3(net326),
.S0(net730),
.S1(net731),
.X(net635)
);

sky130_fd_sc_hd__sdfstp_4 merge740(
.D(net199),
.SCD(net320),
.SCE(net197),
.SET_B(net316),
.CLK(clk),
.Q(net636)
);

sky130_fd_sc_hd__dfxbp_1 s741(
.D(net56),
.CLK(clk),
.Q(out59),
.Q_N(net637)
);

sky130_fd_sc_hd__dfxbp_2 s742(
.D(net60),
.CLK(clk),
.Q(out38),
.Q_N(net638)
);

sky130_fd_sc_hd__dfxtp_1 s743(
.D(net103),
.CLK(clk),
.Q(net639)
);

sky130_fd_sc_hd__dfxtp_2 s744(
.D(net105),
.CLK(clk),
.Q(net640)
);

sky130_fd_sc_hd__dfxtp_4 s745(
.D(net126),
.CLK(clk),
.Q(net641)
);

sky130_fd_sc_hd__dlclkp_1 s746(
.GATE(net129),
.CLK(clk),
.GCLK(net642)
);

sky130_fd_sc_hd__dlclkp_2 s747(
.GATE(net131),
.CLK(clk),
.GCLK(net643)
);

sky130_fd_sc_hd__dlclkp_4 s748(
.GATE(net177),
.CLK(clk),
.GCLK(out12)
);

sky130_fd_sc_hd__dlxbn_1 s749(
.D(net216),
.GATE_N(clk),
.Q(net645),
.Q_N(net644)
);

sky130_fd_sc_hd__dlxbn_2 s750(
.D(net223),
.GATE_N(clk),
.Q(out23),
.Q_N(net646)
);

sky130_fd_sc_hd__dlxbp_1 s751(
.D(net224),
.GATE(clk),
.Q(net648),
.Q_N(net647)
);

sky130_fd_sc_hd__dlxtn_1 s752(
.D(net242),
.GATE_N(clk),
.Q(out17)
);

sky130_fd_sc_hd__dlxtn_2 s753(
.D(net243),
.GATE_N(clk),
.Q(net649)
);

sky130_fd_sc_hd__dlxtn_4 s754(
.D(net263),
.GATE_N(clk),
.Q(net650)
);

sky130_fd_sc_hd__dlxtp_1 s755(
.D(net272),
.GATE(clk),
.Q(out14)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s756(
.D(net273),
.SLEEP_B(clk),
.Q(net651)
);

sky130_fd_sc_hd__dfxbp_1 s757(
.D(net292),
.CLK(clk),
.Q(out36),
.Q_N(net652)
);

sky130_fd_sc_hd__dfxbp_2 s758(
.D(net293),
.CLK(clk),
.Q(out50),
.Q_N(net653)
);

sky130_fd_sc_hd__dfxtp_1 s759(
.D(net294),
.CLK(clk),
.Q(out7)
);

sky130_fd_sc_hd__dfxtp_2 s760(
.D(net295),
.CLK(clk),
.Q(out49)
);

sky130_fd_sc_hd__dfxtp_4 s761(
.D(net296),
.CLK(clk),
.Q(out58)
);

sky130_fd_sc_hd__dlclkp_1 s762(
.GATE(net297),
.CLK(clk),
.GCLK(out53)
);

sky130_fd_sc_hd__dlclkp_2 s763(
.GATE(net368),
.CLK(clk),
.GCLK(out28)
);

sky130_fd_sc_hd__dlclkp_4 s764(
.GATE(net382),
.CLK(clk),
.GCLK(net654)
);

sky130_fd_sc_hd__dlxbn_1 s765(
.D(net383),
.GATE_N(clk),
.Q(net656),
.Q_N(net655)
);

sky130_fd_sc_hd__dlxbn_2 s766(
.D(net386),
.GATE_N(clk),
.Q(net658),
.Q_N(net657)
);

sky130_fd_sc_hd__dlxbp_1 s767(
.D(net387),
.GATE(clk),
.Q(net660),
.Q_N(net659)
);

sky130_fd_sc_hd__dlxtn_1 s768(
.D(net389),
.GATE_N(clk),
.Q(net661)
);

sky130_fd_sc_hd__dlxtn_2 s769(
.D(net390),
.GATE_N(clk),
.Q(net662)
);

sky130_fd_sc_hd__dlxtn_4 s770(
.D(net391),
.GATE_N(clk),
.Q(net663)
);

sky130_fd_sc_hd__dlxtp_1 s771(
.D(net392),
.GATE(clk),
.Q(net664)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s772(
.D(net400),
.SLEEP_B(clk),
.Q(net665)
);

sky130_fd_sc_hd__dfxbp_1 s773(
.D(net402),
.CLK(clk),
.Q(out16),
.Q_N(net666)
);

sky130_fd_sc_hd__dfxbp_2 s774(
.D(net403),
.CLK(clk),
.Q(net667)
);

sky130_fd_sc_hd__dfxtp_1 s775(
.D(net404),
.CLK(clk),
.Q(out41)
);

sky130_fd_sc_hd__dfxtp_2 s776(
.D(net405),
.CLK(clk),
.Q(net668)
);

sky130_fd_sc_hd__dfxtp_4 s777(
.D(net427),
.CLK(clk),
.Q(net669)
);

sky130_fd_sc_hd__dlclkp_1 s778(
.GATE(net431),
.CLK(clk),
.GCLK(net670)
);

sky130_fd_sc_hd__dlclkp_2 s779(
.GATE(net464),
.CLK(clk),
.GCLK(net671)
);

sky130_fd_sc_hd__dlclkp_4 s780(
.GATE(net473),
.CLK(clk),
.GCLK(net672)
);

sky130_fd_sc_hd__dlxbn_1 s781(
.D(net475),
.GATE_N(clk),
.Q(net673)
);

sky130_fd_sc_hd__dlxbn_2 s782(
.D(net477),
.GATE_N(clk),
.Q(net675),
.Q_N(net674)
);

sky130_fd_sc_hd__dlxbp_1 s783(
.D(net478),
.GATE(clk),
.Q(net677),
.Q_N(net676)
);

sky130_fd_sc_hd__dlxtn_1 s784(
.D(net480),
.GATE_N(clk),
.Q(net678)
);

sky130_fd_sc_hd__dlxtn_2 s785(
.D(net481),
.GATE_N(clk),
.Q(net679)
);

sky130_fd_sc_hd__dlxtn_4 s786(
.D(net488),
.GATE_N(clk),
.Q(net680)
);

sky130_fd_sc_hd__dlxtp_1 s787(
.D(net495),
.GATE(clk),
.Q(net681)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s788(
.D(net497),
.SLEEP_B(clk),
.Q(net682)
);

sky130_fd_sc_hd__dfxbp_1 s789(
.D(net499),
.CLK(clk),
.Q(net684),
.Q_N(net683)
);

sky130_fd_sc_hd__dfxbp_2 s790(
.D(net500),
.CLK(clk),
.Q(net686),
.Q_N(net685)
);

sky130_fd_sc_hd__dfxtp_1 s791(
.D(net502),
.CLK(clk),
.Q(net687)
);

sky130_fd_sc_hd__dfxtp_2 s792(
.D(net507),
.CLK(clk),
.Q(net688)
);

sky130_fd_sc_hd__dfxtp_4 s793(
.D(net509),
.CLK(clk),
.Q(out20)
);

sky130_fd_sc_hd__dlclkp_1 s794(
.GATE(net510),
.CLK(clk),
.GCLK(net689)
);

sky130_fd_sc_hd__dlclkp_2 s795(
.GATE(net515),
.CLK(clk),
.GCLK(net690)
);

sky130_fd_sc_hd__dlclkp_4 s796(
.GATE(net516),
.CLK(clk),
.GCLK(net691)
);

sky130_fd_sc_hd__dlxbn_1 s797(
.D(net518),
.GATE_N(clk),
.Q(net693),
.Q_N(net692)
);

sky130_fd_sc_hd__dlxbn_2 s798(
.D(net519),
.GATE_N(clk),
.Q(out11),
.Q_N(net694)
);

sky130_fd_sc_hd__dlxbp_1 s799(
.D(net520),
.GATE(clk),
.Q(net696),
.Q_N(net695)
);

sky130_fd_sc_hd__dlxtn_1 s800(
.D(net521),
.GATE_N(clk),
.Q(net697)
);

sky130_fd_sc_hd__dlxtn_2 s801(
.D(net523),
.GATE_N(clk),
.Q(net698)
);

sky130_fd_sc_hd__dlxtn_4 s802(
.D(net544),
.GATE_N(clk),
.Q(out3)
);

sky130_fd_sc_hd__dlxtp_1 s803(
.D(net545),
.GATE(clk),
.Q(net699)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s804(
.D(net556),
.SLEEP_B(clk),
.Q(net700)
);

sky130_fd_sc_hd__dfxbp_1 s805(
.D(net571),
.CLK(clk),
.Q(net701)
);

sky130_fd_sc_hd__dfxbp_2 s806(
.D(net574),
.CLK(clk),
.Q(net702)
);

sky130_fd_sc_hd__dfxtp_1 s807(
.D(net579),
.CLK(clk),
.Q(net703)
);

sky130_fd_sc_hd__dfxtp_2 s808(
.D(net584),
.CLK(clk),
.Q(net704)
);

sky130_fd_sc_hd__dfxtp_4 s809(
.D(net588),
.CLK(clk),
.Q(net705)
);

sky130_fd_sc_hd__dlclkp_1 s810(
.GATE(net591),
.CLK(clk),
.GCLK(net706)
);

sky130_fd_sc_hd__dlclkp_2 s811(
.GATE(net598),
.CLK(clk),
.GCLK(net707)
);

sky130_fd_sc_hd__dlclkp_4 s812(
.GATE(net599),
.CLK(clk),
.GCLK(net708)
);

sky130_fd_sc_hd__dlxbn_1 s813(
.D(net601),
.GATE_N(clk),
.Q(net710),
.Q_N(net709)
);

sky130_fd_sc_hd__dlxbn_2 s814(
.D(net603),
.GATE_N(clk),
.Q(net712),
.Q_N(net711)
);

sky130_fd_sc_hd__dlxbp_1 s815(
.D(net605),
.GATE(clk),
.Q(net714),
.Q_N(net713)
);

sky130_fd_sc_hd__dlxtn_1 s816(
.D(net608),
.GATE_N(clk),
.Q(net715)
);

sky130_fd_sc_hd__dlxtn_2 s817(
.D(net611),
.GATE_N(clk),
.Q(net716)
);

sky130_fd_sc_hd__dlxtn_4 s818(
.D(net612),
.GATE_N(clk),
.Q(net717)
);

sky130_fd_sc_hd__dlxtp_1 s819(
.D(net613),
.GATE(clk),
.Q(net718)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s820(
.D(net616),
.SLEEP_B(clk),
.Q(net719)
);

sky130_fd_sc_hd__dfxbp_1 s821(
.D(net617),
.CLK(clk),
.Q(net720)
);

sky130_fd_sc_hd__dfxbp_2 s822(
.D(net621),
.CLK(clk),
.Q(net721)
);

sky130_fd_sc_hd__dfxtp_1 s823(
.D(net623),
.CLK(clk),
.Q(net722)
);

sky130_fd_sc_hd__dfxtp_2 s824(
.D(net624),
.CLK(clk),
.Q(net723)
);

sky130_fd_sc_hd__dfxtp_4 s825(
.D(net625),
.CLK(clk),
.Q(net724)
);

sky130_fd_sc_hd__dlclkp_1 s826(
.GATE(net626),
.CLK(clk),
.GCLK(net725)
);

sky130_fd_sc_hd__dlclkp_2 s827(
.GATE(net627),
.CLK(clk),
.GCLK(net726)
);

sky130_fd_sc_hd__dlclkp_4 s828(
.GATE(net629),
.CLK(clk),
.GCLK(net727)
);

sky130_fd_sc_hd__dlxbn_1 s829(
.D(net630),
.GATE_N(clk),
.Q(net728)
);

sky130_fd_sc_hd__dlxbn_2 s830(
.D(net632),
.GATE_N(clk),
.Q(net729)
);

sky130_fd_sc_hd__dlxbp_1 s831(
.D(net633),
.GATE(clk),
.Q(net730)
);

sky130_fd_sc_hd__dlxtn_1 s832(
.D(net634),
.GATE_N(clk),
.Q(net731)
);

sky130_fd_sc_hd__dlxtn_2 s833(
.D(net635),
.GATE_N(clk)
);


endmodule
