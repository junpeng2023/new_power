module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net995;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire clknet_0_clk;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net978;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net987;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net996;
 wire net997;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net814;
 wire clknet_1_0__leaf_net814;
 wire clknet_1_1__leaf_net814;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net599;
 wire clknet_1_0__leaf_net599;
 wire clknet_1_1__leaf_net599;
 wire clknet_0_net598;
 wire clknet_1_0__leaf_net598;
 wire clknet_1_1__leaf_net598;
 wire clknet_0_net813;
 wire clknet_1_0__leaf_net813;
 wire clknet_1_1__leaf_net813;
 wire clknet_0_net812;
 wire clknet_1_0__leaf_net812;
 wire clknet_1_1__leaf_net812;
 wire clknet_0_net940;
 wire clknet_1_0__leaf_net940;
 wire clknet_1_1__leaf_net940;
 wire clknet_0_net638;
 wire clknet_1_0__leaf_net638;
 wire clknet_1_1__leaf_net638;
 wire clknet_0_net643;
 wire clknet_1_0__leaf_net643;
 wire clknet_1_1__leaf_net643;
 wire clknet_0_net904;
 wire clknet_1_0__leaf_net904;
 wire clknet_1_1__leaf_net904;
 wire clknet_0_net795;
 wire clknet_1_0__leaf_net795;
 wire clknet_1_1__leaf_net795;
 wire clknet_0_net901;
 wire clknet_1_0__leaf_net901;
 wire clknet_1_1__leaf_net901;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net182;
 wire clknet_1_0__leaf_net182;
 wire clknet_1_1__leaf_net182;
 wire clknet_0_net776;
 wire clknet_1_0__leaf_net776;
 wire clknet_1_1__leaf_net776;
 wire clknet_0_net135;
 wire clknet_1_0__leaf_net135;
 wire clknet_1_1__leaf_net135;
 wire clknet_0_net894;
 wire clknet_1_0__leaf_net894;
 wire clknet_1_1__leaf_net894;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net933;
 wire clknet_1_0__leaf_net933;
 wire clknet_1_1__leaf_net933;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net292;
 wire clknet_1_0__leaf_net292;
 wire clknet_1_1__leaf_net292;
 wire clknet_0_net286;
 wire clknet_1_0__leaf_net286;
 wire clknet_1_1__leaf_net286;
 wire clknet_0_net748;
 wire clknet_1_0__leaf_net748;
 wire clknet_1_1__leaf_net748;
 wire clknet_0_net414;
 wire clknet_1_0__leaf_net414;
 wire clknet_1_1__leaf_net414;
 wire clknet_0_net423;
 wire clknet_1_0__leaf_net423;
 wire clknet_1_1__leaf_net423;
 wire clknet_0_net905;
 wire clknet_1_0__leaf_net905;
 wire clknet_1_1__leaf_net905;
 wire clknet_0_net937;
 wire clknet_1_0__leaf_net937;
 wire clknet_1_1__leaf_net937;
 wire clknet_0_net777;
 wire clknet_1_0__leaf_net777;
 wire clknet_1_1__leaf_net777;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net291;
 wire clknet_1_0__leaf_net291;
 wire clknet_1_1__leaf_net291;
 wire clknet_0_net747;
 wire clknet_1_0__leaf_net747;
 wire clknet_1_1__leaf_net747;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net407;
 wire clknet_1_0__leaf_net407;
 wire clknet_1_1__leaf_net407;
 wire clknet_0_net394;
 wire clknet_1_0__leaf_net394;
 wire clknet_1_1__leaf_net394;
 wire clknet_0_net276;
 wire clknet_1_0__leaf_net276;
 wire clknet_1_1__leaf_net276;
 wire clknet_0_net148;
 wire clknet_1_0__leaf_net148;
 wire clknet_1_1__leaf_net148;
 wire clknet_0_net145;
 wire clknet_1_0__leaf_net145;
 wire clknet_1_1__leaf_net145;
 wire clknet_0_net146;
 wire clknet_1_0__leaf_net146;
 wire clknet_1_1__leaf_net146;
 wire clknet_0_net140;
 wire clknet_1_0__leaf_net140;
 wire clknet_1_1__leaf_net140;
 wire clknet_0_net153;
 wire clknet_1_0__leaf_net153;
 wire clknet_1_1__leaf_net153;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire clknet_0_net169;
 wire clknet_1_0__leaf_net169;
 wire clknet_1_1__leaf_net169;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net921;
 wire clknet_1_0__leaf_net921;
 wire clknet_1_1__leaf_net921;
 wire clknet_0_net143;
 wire clknet_1_0__leaf_net143;
 wire clknet_1_1__leaf_net143;
 wire clknet_0_net395;
 wire clknet_1_0__leaf_net395;
 wire clknet_1_1__leaf_net395;
 wire clknet_0_net939;
 wire clknet_1_0__leaf_net939;
 wire clknet_1_1__leaf_net939;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net152;
 wire clknet_1_0__leaf_net152;
 wire clknet_1_1__leaf_net152;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net136;
 wire clknet_1_0__leaf_net136;
 wire clknet_1_1__leaf_net136;
 wire clknet_0_net406;
 wire clknet_1_0__leaf_net406;
 wire clknet_1_1__leaf_net406;
 wire clknet_0_net516;
 wire clknet_1_0__leaf_net516;
 wire clknet_1_1__leaf_net516;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net910;
 wire clknet_1_0__leaf_net910;
 wire clknet_1_1__leaf_net910;
 wire clknet_0_net920;
 wire clknet_1_0__leaf_net920;
 wire clknet_1_1__leaf_net920;
 wire clknet_0_net306;
 wire clknet_1_0__leaf_net306;
 wire clknet_1_1__leaf_net306;
 wire clknet_0_net425;
 wire clknet_1_0__leaf_net425;
 wire clknet_1_1__leaf_net425;
 wire clknet_0_net794;
 wire clknet_1_0__leaf_net794;
 wire clknet_1_1__leaf_net794;
 wire clknet_0_net564;
 wire clknet_1_0__leaf_net564;
 wire clknet_1_1__leaf_net564;
 wire clknet_0_net584;
 wire clknet_1_0__leaf_net584;
 wire clknet_1_1__leaf_net584;
 wire clknet_0_net575;
 wire clknet_1_0__leaf_net575;
 wire clknet_1_1__leaf_net575;
 wire clknet_0_net570;
 wire clknet_1_0__leaf_net570;
 wire clknet_1_1__leaf_net570;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net563;
 wire clknet_0_net387;
 wire clknet_1_0__leaf_net387;
 wire clknet_1_1__leaf_net387;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net371;
 wire clknet_1_0__leaf_net371;
 wire clknet_1_1__leaf_net371;
 wire clknet_0_net366;
 wire clknet_1_0__leaf_net366;
 wire clknet_1_1__leaf_net366;
 wire clknet_0_net527;
 wire clknet_1_0__leaf_net527;
 wire clknet_1_1__leaf_net527;
 wire clknet_0_net917;
 wire clknet_1_0__leaf_net917;
 wire clknet_1_1__leaf_net917;
 wire clknet_0_net382;
 wire clknet_1_0__leaf_net382;
 wire clknet_1_1__leaf_net382;
 wire clknet_0_net363;
 wire clknet_1_0__leaf_net363;
 wire clknet_1_1__leaf_net363;
 wire clknet_0_net460;
 wire clknet_1_0__leaf_net460;
 wire clknet_1_1__leaf_net460;
 wire clknet_0_net452;
 wire clknet_1_0__leaf_net452;
 wire clknet_1_1__leaf_net452;
 wire clknet_0_net439;
 wire clknet_1_0__leaf_net439;
 wire clknet_1_1__leaf_net439;
 wire clknet_0_net552;
 wire clknet_1_0__leaf_net552;
 wire clknet_1_1__leaf_net552;
 wire clknet_0_net440;
 wire clknet_1_0__leaf_net440;
 wire clknet_1_1__leaf_net440;
 wire clknet_0_net478;
 wire clknet_1_0__leaf_net478;
 wire clknet_1_1__leaf_net478;
 wire clknet_0_net477;
 wire clknet_1_0__leaf_net477;
 wire clknet_1_1__leaf_net477;
 wire clknet_0_net472;
 wire clknet_1_0__leaf_net472;
 wire clknet_1_1__leaf_net472;
 wire clknet_0_net447;
 wire clknet_1_0__leaf_net447;
 wire clknet_1_1__leaf_net447;
 wire clknet_0_net442;
 wire clknet_1_0__leaf_net442;
 wire clknet_1_1__leaf_net442;
 wire clknet_0_net445;
 wire clknet_1_0__leaf_net445;
 wire clknet_1_1__leaf_net445;
 wire clknet_0_net438;
 wire clknet_1_0__leaf_net438;
 wire clknet_1_1__leaf_net438;
 wire clknet_0_net899;
 wire clknet_1_0__leaf_net899;
 wire clknet_1_1__leaf_net899;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net379;
 wire clknet_1_0__leaf_net379;
 wire clknet_1_1__leaf_net379;
 wire clknet_0_net373;
 wire clknet_1_0__leaf_net373;
 wire clknet_1_1__leaf_net373;
 wire clknet_0_net254;
 wire clknet_1_0__leaf_net254;
 wire clknet_1_1__leaf_net254;
 wire net131;
 wire net227;
 wire net436;
 wire net912;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;

 sky130_fd_sc_hd__nand2b_1 c100 (.A_N(net29),
    .B(net958),
    .Y(net36));
 sky130_fd_sc_hd__nor2_4 c101 (.A(net18),
    .B(net958),
    .Y(net37));
 sky130_fd_sc_hd__nor2b_2 c102 (.A(net923),
    .B_N(net32),
    .Y(net38));
 sky130_fd_sc_hd__o2111ai_4 c103 (.A1(net14),
    .A2(net29),
    .B1(net957),
    .C1(net828),
    .D1(net31),
    .Y(net932));
 sky130_fd_sc_hd__and2b_1 c104 (.A_N(net36),
    .B(net18),
    .X(net39));
 sky130_fd_sc_hd__a2111oi_1 c105 (.A1(net959),
    .A2(net29),
    .B1(net37),
    .C1(net18),
    .D1(net35),
    .Y(net40));
 sky130_fd_sc_hd__or4bb_1 c106 (.A(net39),
    .B(net959),
    .C_N(net40),
    .D_N(net35),
    .X(net41));
 sky130_fd_sc_hd__a2111o_4 c107 (.A1(net28),
    .A2(net37),
    .B1(net932),
    .C1(net38),
    .D1(net32),
    .X(net42));
 sky130_fd_sc_hd__nand2_2 c108 (.A(net41),
    .B(net37),
    .Y(net43));
 sky130_fd_sc_hd__nor2_4 c109 (.A(net956),
    .B(net932),
    .Y(net931));
 sky130_fd_sc_hd__nor2_1 c110 (.A(net841),
    .B(net21),
    .Y(net44));
 sky130_fd_sc_hd__and2_2 c111 (.A(net828),
    .B(net835),
    .X(net45));
 sky130_fd_sc_hd__nor2b_1 c112 (.A(net28),
    .B_N(net16),
    .Y(net46));
 sky130_fd_sc_hd__nand2_2 c113 (.A(net861),
    .B(net44),
    .Y(net47));
 sky130_fd_sc_hd__and2b_1 c114 (.A_N(net32),
    .B(net34),
    .X(net48));
 sky130_fd_sc_hd__and2b_2 c115 (.A_N(net16),
    .B(net28),
    .X(net908));
 sky130_fd_sc_hd__or2_2 c116 (.A(net870),
    .B(net972),
    .X(net49));
 sky130_fd_sc_hd__nor2_1 c117 (.A(net44),
    .B(net26),
    .Y(net50));
 sky130_fd_sc_hd__and2_2 c118 (.A(net47),
    .B(net49),
    .X(net891));
 sky130_fd_sc_hd__nor3b_1 c119 (.A(net50),
    .B(net44),
    .C_N(net48),
    .Y(net51));
 sky130_fd_sc_hd__and2_1 c120 (.A(net891),
    .B(net21),
    .X(net52));
 sky130_fd_sc_hd__or4bb_1 c121 (.A(net972),
    .B(net873),
    .C_N(net52),
    .D_N(net870),
    .X(net53));
 sky130_fd_sc_hd__and2_0 c122 (.A(net52),
    .B(net891),
    .X(net54));
 sky130_fd_sc_hd__and2b_2 c123 (.A_N(net26),
    .B(net49),
    .X(net55));
 sky130_fd_sc_hd__o2111ai_1 c124 (.A1(net51),
    .A2(net908),
    .B1(net53),
    .C1(net891),
    .D1(net45),
    .Y(net56));
 sky130_fd_sc_hd__mux4_2 c125 (.A0(net53),
    .A1(net862),
    .A2(net46),
    .A3(net891),
    .S0(net844),
    .S1(net55),
    .X(net57));
 sky130_fd_sc_hd__or4bb_1 c126 (.A(net21),
    .B(net52),
    .C_N(net34),
    .D_N(net49),
    .X(net58));
 sky130_fd_sc_hd__and3b_4 c127 (.A_N(net54),
    .B(net908),
    .C(net50),
    .X(net925));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net48),
    .A1(net54),
    .A2(net55),
    .A3(net925),
    .S0(net58),
    .S1(net49),
    .X(net59));
 sky130_fd_sc_hd__and2b_1 c129 (.A_N(net53),
    .B(net925),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net58),
    .A1(net60),
    .A2(net56),
    .A3(net925),
    .S0(net891),
    .S1(net59),
    .X(net61));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net57),
    .A1(net59),
    .A2(net51),
    .A3(net925),
    .S0(net55),
    .S1(net58),
    .X(net62));
 sky130_fd_sc_hd__nand2b_4 c132 (.A_N(net830),
    .B(net836),
    .Y(net63));
 sky130_fd_sc_hd__nor3_2 c133 (.A(net63),
    .B(net883),
    .C(net884),
    .Y(net64));
 sky130_fd_sc_hd__nor2b_4 c134 (.A(net64),
    .B_N(net824),
    .Y(net65));
 sky130_fd_sc_hd__or2_1 c135 (.A(net884),
    .B(net64),
    .X(net66));
 sky130_fd_sc_hd__nand2b_4 c136 (.A_N(net64),
    .B(net65),
    .Y(net67));
 sky130_fd_sc_hd__nor3b_4 c137 (.A(net834),
    .B(net827),
    .C_N(net825),
    .Y(net68));
 sky130_fd_sc_hd__or2b_4 c138 (.A(net67),
    .B_N(net825),
    .X(net69));
 sky130_fd_sc_hd__nor2b_1 c139 (.A(net880),
    .B_N(net66),
    .Y(net70));
 sky130_fd_sc_hd__and2_4 c140 (.A(net69),
    .B(net68),
    .X(net71));
 sky130_fd_sc_hd__and2b_4 c141 (.A_N(net883),
    .B(net836),
    .X(net72));
 sky130_fd_sc_hd__mux4_2 c142 (.A0(net70),
    .A1(net71),
    .A2(net834),
    .A3(net72),
    .S0(net65),
    .S1(net824),
    .X(net73));
 sky130_fd_sc_hd__nor2b_2 c143 (.A(net68),
    .B_N(net63),
    .Y(net74));
 sky130_fd_sc_hd__and3_2 c144 (.A(net74),
    .B(net68),
    .C(net72),
    .X(net75));
 sky130_fd_sc_hd__and2_2 c145 (.A(net73),
    .B(net70),
    .X(net76));
 sky130_fd_sc_hd__nand3b_4 c146 (.A_N(net75),
    .B(net73),
    .C(net830),
    .Y(net77));
 sky130_fd_sc_hd__and2_4 c147 (.A(net77),
    .B(net824),
    .X(net78));
 sky130_fd_sc_hd__or4bb_4 c148 (.A(net77),
    .B(net66),
    .C_N(net68),
    .D_N(net71),
    .X(net79));
 sky130_fd_sc_hd__mux4_2 c149 (.A0(net825),
    .A1(net73),
    .A2(net824),
    .A3(net68),
    .S0(net885),
    .S1(net880),
    .X(net80));
 sky130_fd_sc_hd__or3_2 c150 (.A(net227),
    .B(net869),
    .C(net76),
    .X(net81));
 sky130_fd_sc_hd__nand3_4 c151 (.A(net76),
    .B(net81),
    .C(net63),
    .Y(net82));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net63),
    .A1(net80),
    .A2(net847),
    .A3(net74),
    .S0(net76),
    .S1(net82),
    .X(net900));
 sky130_fd_sc_hd__nor3b_4 c153 (.A(net79),
    .B(net80),
    .C_N(net69),
    .Y(net83));
 sky130_fd_sc_hd__nor3b_2 c154 (.A(net869),
    .B(net832),
    .C_N(net847),
    .Y(net84));
 sky130_fd_sc_hd__nand3b_4 c155 (.A_N(net81),
    .B(net68),
    .C(net836),
    .Y(net85));
 sky130_fd_sc_hd__or2b_1 c156 (.A(net854),
    .B_N(net81),
    .X(net86));
 sky130_fd_sc_hd__nor3b_1 c157 (.A(net843),
    .B(net85),
    .C_N(net80),
    .Y(net87));
 sky130_fd_sc_hd__nor3b_2 c158 (.A(net832),
    .B(net859),
    .C_N(net851),
    .Y(net88));
 sky130_fd_sc_hd__and2_1 c159 (.A(net73),
    .B(net848),
    .X(net89));
 sky130_fd_sc_hd__nor3b_2 c160 (.A(net80),
    .B(net855),
    .C_N(net859),
    .Y(net90));
 sky130_fd_sc_hd__or2_1 c161 (.A(net855),
    .B(net68),
    .X(net91));
 sky130_fd_sc_hd__nand2_1 c162 (.A(net831),
    .B(net83),
    .Y(net92));
 sky130_fd_sc_hd__or2b_2 c163 (.A(net860),
    .B_N(net844),
    .X(net93));
 sky130_fd_sc_hd__nor2b_1 c164 (.A(net853),
    .B_N(net85),
    .Y(net94));
 sky130_fd_sc_hd__a2111o_2 c165 (.A1(net837),
    .A2(net94),
    .B1(net86),
    .C1(net227),
    .D1(net67),
    .X(net95));
 sky130_fd_sc_hd__nand3b_2 c166 (.A_N(net829),
    .B(net859),
    .C(net973),
    .Y(net96));
 sky130_fd_sc_hd__nor3b_4 c167 (.A(net96),
    .B(net973),
    .C_N(net89),
    .Y(net97));
 sky130_fd_sc_hd__and2_1 c168 (.A(net86),
    .B(net65),
    .X(net98));
 sky130_fd_sc_hd__or4bb_1 c169 (.A(net89),
    .B(net79),
    .C_N(net97),
    .D_N(net973),
    .X(net99));
 sky130_fd_sc_hd__and3_1 c170 (.A(net98),
    .B(net99),
    .C(net86),
    .X(net100));
 sky130_fd_sc_hd__and3b_2 c171 (.A_N(net858),
    .B(net96),
    .C(net98),
    .X(net918));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net92),
    .A1(net100),
    .A2(net85),
    .A3(net88),
    .S0(net852),
    .S1(net857),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net94),
    .A1(net862),
    .A2(net973),
    .A3(net101),
    .S0(net79),
    .S1(net951),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net68),
    .A1(net101),
    .A2(net102),
    .A3(net85),
    .S0(net846),
    .S1(net86),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net100),
    .A1(net91),
    .A2(net859),
    .A3(net102),
    .S0(net101),
    .X(net104));
 sky130_fd_sc_hd__nor3b_4 c176 (.A(net881),
    .B(net874),
    .C_N(net870),
    .Y(net105));
 sky130_fd_sc_hd__or3_4 c177 (.A(net96),
    .B(net85),
    .C(net848),
    .X(net106));
 sky130_fd_sc_hd__or4bb_1 c178 (.A(net92),
    .B(net881),
    .C_N(net84),
    .D_N(net900),
    .X(net107));
 sky130_fd_sc_hd__or4bb_4 c179 (.A(net852),
    .B(net96),
    .C_N(net847),
    .D_N(net878),
    .X(net108));
 sky130_fd_sc_hd__and3_1 c180 (.A(net105),
    .B(net106),
    .C(net689),
    .X(net109));
 sky130_fd_sc_hd__or3_1 c181 (.A(net82),
    .B(net109),
    .C(net689),
    .X(net110));
 sky130_fd_sc_hd__nand3b_1 c182 (.A_N(net882),
    .B(net82),
    .C(net87),
    .Y(net111));
 sky130_fd_sc_hd__and3_1 c183 (.A(net848),
    .B(net873),
    .C(net110),
    .X(net112));
 sky130_fd_sc_hd__nor3_1 c184 (.A(net107),
    .B(net108),
    .C(net105),
    .Y(net113));
 sky130_fd_sc_hd__or4bb_1 c185 (.A(net108),
    .B(net852),
    .C_N(net113),
    .D_N(net951),
    .X(net114));
 sky130_fd_sc_hd__or3b_1 c186 (.A(net848),
    .B(net877),
    .C_N(net108),
    .X(net115));
 sky130_fd_sc_hd__or4bb_2 c187 (.A(net109),
    .B(net111),
    .C_N(net862),
    .D_N(net689),
    .X(net116));
 sky130_fd_sc_hd__inv_2 c188 (.A(net743),
    .Y(net117));
 sky130_fd_sc_hd__mux4_1 c189 (.A0(net87),
    .A1(net112),
    .A2(net2),
    .A3(net115),
    .S0(net969),
    .S1(net864),
    .X(net118));
 sky130_fd_sc_hd__or4bb_1 c190 (.A(net115),
    .B(net116),
    .C_N(net850),
    .D_N(net742),
    .X(net119));
 sky130_fd_sc_hd__o2111a_2 c191 (.A1(net97),
    .A2(net115),
    .B1(net969),
    .C1(net105),
    .D1(net108),
    .X(net120));
 sky130_fd_sc_hd__or4bb_1 c192 (.A(net113),
    .B(net107),
    .C_N(net108),
    .D_N(net742),
    .X(net121));
 sky130_fd_sc_hd__sdfrbp_2 c193 (.CLK(clknet_4_2_0_clk),
    .D(net121),
    .RESET_B(net109),
    .SCD(net75),
    .SCE(net969),
    .Q(net123),
    .Q_N(net122));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net110),
    .A1(net877),
    .A2(net879),
    .A3(net876),
    .S0(net108),
    .S1(net742),
    .X(net124));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net109),
    .A1(net108),
    .A2(net969),
    .A3(net124),
    .S0(net122),
    .S1(net743),
    .X(net125));
 sky130_fd_sc_hd__mux4_2 c196 (.A0(net116),
    .A1(net873),
    .A2(net969),
    .A3(net122),
    .S0(net742),
    .S1(net788),
    .X(net126));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net124),
    .A1(net123),
    .A2(net97),
    .A3(net969),
    .S0(net742),
    .S1(net787),
    .X(net127));
 sky130_fd_sc_hd__nand3_4 c198 (.A(net866),
    .B(net949),
    .C(net23),
    .Y(net128));
 sky130_fd_sc_hd__nand2b_1 c199 (.A_N(net1),
    .B(net857),
    .Y(net129));
 sky130_fd_sc_hd__clkbuf_1 c200 (.A(net704),
    .X(net130));
 sky130_fd_sc_hd__clkinv_1 c301_21 (.A(clknet_1_0__leaf_net776),
    .Y(net995));
 sky130_fd_sc_hd__or3b_1 c202 (.A(net1024),
    .B(net120),
    .C_N(net951),
    .X(net132));
 sky130_fd_sc_hd__clkinv_8 c203 (.A(net734),
    .Y(net133));
 sky130_fd_sc_hd__inv_4 c204 (.A(net704),
    .Y(net134));
 sky130_fd_sc_hd__nand3_4 c205 (.A(net994),
    .B(net974),
    .C(net133),
    .Y(net135));
 sky130_fd_sc_hd__a2111o_2 c206 (.A1(net864),
    .A2(clknet_1_0__leaf_net135),
    .B1(net227),
    .C1(net134),
    .D1(net961),
    .X(net136));
 sky130_fd_sc_hd__a2111oi_2 c207 (.A1(net83),
    .A2(net8),
    .B1(net969),
    .C1(net862),
    .D1(net23),
    .Y(net137));
 sky130_fd_sc_hd__clkbuf_4 c208 (.A(net704),
    .X(net138));
 sky130_fd_sc_hd__or3_1 c209 (.A(net849),
    .B(net970),
    .C(net133),
    .X(net139));
 sky130_fd_sc_hd__mux4_2 c210 (.A0(clknet_1_0__leaf_net136),
    .A1(net23),
    .A2(net88),
    .A3(net993),
    .S0(net138),
    .S1(clknet_1_1__leaf_net135),
    .X(net140));
 sky130_fd_sc_hd__a2111oi_1 c211 (.A1(net139),
    .A2(net83),
    .B1(net69),
    .C1(net961),
    .D1(net787),
    .Y(net141));
 sky130_fd_sc_hd__nand3_1 c212 (.A(net954),
    .B(net120),
    .C(clknet_1_1__leaf_net140),
    .Y(net142));
 sky130_fd_sc_hd__a2111o_2 c213 (.A1(net137),
    .A2(net139),
    .B1(net1004),
    .C1(clknet_1_0__leaf_net142),
    .D1(clknet_1_0__leaf_net135),
    .X(net894));
 sky130_fd_sc_hd__or3_4 c214 (.A(clknet_1_0__leaf_net140),
    .B(net955),
    .C(net134),
    .X(net143));
 sky130_fd_sc_hd__mux4_4 c215 (.A0(net8),
    .A1(clknet_1_0__leaf_net143),
    .A2(net91),
    .A3(net949),
    .S0(net1),
    .S1(net128),
    .X(net144));
 sky130_fd_sc_hd__mux4_2 c216 (.A0(clknet_1_0__leaf_net142),
    .A1(clknet_1_1__leaf_net136),
    .A2(net138),
    .A3(clknet_1_0__leaf_net140),
    .S0(clknet_1_0__leaf_net894),
    .S1(net734),
    .X(net145));
 sky130_fd_sc_hd__mux4_2 c217 (.A0(net874),
    .A1(net133),
    .A2(clknet_1_0__leaf_net145),
    .A3(net23),
    .S0(net138),
    .S1(net734),
    .X(net146));
 sky130_fd_sc_hd__inv_4 c218 (.A(net704),
    .Y(net147));
 sky130_fd_sc_hd__a2111o_1 c219 (.A1(clknet_1_1__leaf_net145),
    .A2(net147),
    .B1(net840),
    .C1(net120),
    .D1(clknet_1_0__leaf_net894),
    .X(net148));
 sky130_fd_sc_hd__and2b_1 c220 (.A_N(net132),
    .B(net827),
    .X(net149));
 sky130_fd_sc_hd__nor3_4 c221 (.A(clknet_1_0__leaf_net140),
    .B(net974),
    .C(net957),
    .Y(net921));
 sky130_fd_sc_hd__or2b_2 c222 (.A(net961),
    .B_N(net838),
    .X(net150));
 sky130_fd_sc_hd__nor2b_1 c223 (.A(net130),
    .B_N(net69),
    .Y(net151));
 sky130_fd_sc_hd__o2111a_2 c224 (.A1(clknet_1_1__leaf_net142),
    .A2(net42),
    .B1(net957),
    .C1(net37),
    .D1(net958),
    .X(net152));
 sky130_fd_sc_hd__nor2b_4 c225 (.A(net974),
    .B_N(clknet_1_1__leaf_net140),
    .Y(net153));
 sky130_fd_sc_hd__nand2_4 c226 (.A(net869),
    .B(net23),
    .Y(net154));
 sky130_fd_sc_hd__or3b_1 c227 (.A(net954),
    .B(net154),
    .C_N(net150),
    .X(net155));
 sky130_fd_sc_hd__nand3_2 c228 (.A(clknet_1_0__leaf_net153),
    .B(net931),
    .C(net43),
    .Y(net156));
 sky130_fd_sc_hd__and3b_1 c229 (.A_N(net949),
    .B(net37),
    .C(net155),
    .X(net157));
 sky130_fd_sc_hd__sdfrbp_2 c230 (.CLK(clknet_4_8_0_clk),
    .D(clknet_1_1__leaf_net152),
    .RESET_B(net157),
    .SCD(clknet_1_0__leaf_net156),
    .SCE(net150),
    .Q(net927),
    .Q_N(net158));
 sky130_fd_sc_hd__inv_6 c231 (.A(net741),
    .Y(net159));
 sky130_fd_sc_hd__mux4_2 c232 (.A0(clknet_1_0__leaf_net156),
    .A1(net19),
    .A2(net158),
    .A3(net154),
    .S0(net105),
    .S1(net961),
    .X(net160));
 sky130_fd_sc_hd__o2111ai_1 c233 (.A1(net827),
    .A2(net838),
    .B1(net927),
    .C1(net154),
    .D1(clknet_1_0__leaf_net152),
    .Y(net161));
 sky130_fd_sc_hd__clkinv_8 c234 (.A(net741),
    .Y(net162));
 sky130_fd_sc_hd__sdfrtn_1 c235 (.CLK_N(clknet_4_10_0_clk),
    .D(net159),
    .RESET_B(clknet_1_1__leaf_net161),
    .SCD(net162),
    .SCE(net35),
    .Q(net163));
 sky130_fd_sc_hd__clkbuf_1 c236 (.A(net762),
    .X(net164));
 sky130_fd_sc_hd__sdfrtp_1 c237 (.CLK(clknet_4_8_0_clk),
    .D(net164),
    .RESET_B(net132),
    .SCD(clknet_1_0__leaf_net921),
    .SCE(net149),
    .Q(net165));
 sky130_fd_sc_hd__or4bb_1 c238 (.A(net151),
    .B(net162),
    .C_N(net165),
    .D_N(net159),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net165),
    .A1(clknet_1_1__leaf_net148),
    .A2(net2),
    .A3(net158),
    .S0(net833),
    .S1(net120),
    .X(net167));
 sky130_fd_sc_hd__a2111oi_0 c240 (.A1(net162),
    .A2(net165),
    .B1(clknet_1_0__leaf_net161),
    .C1(clknet_1_1__leaf_net156),
    .D1(net150),
    .Y(net168));
 sky130_fd_sc_hd__o2111ai_2 c241 (.A1(clknet_1_1__leaf_net156),
    .A2(net162),
    .B1(net165),
    .C1(net873),
    .D1(net741),
    .Y(net169));
 sky130_fd_sc_hd__and3b_1 c242 (.A_N(net34),
    .B(net55),
    .C(net958),
    .X(net170));
 sky130_fd_sc_hd__mux4_2 c243 (.A0(clknet_1_0__leaf_net169),
    .A1(net150),
    .A2(net38),
    .A3(net57),
    .S0(net908),
    .S1(net958),
    .X(net171));
 sky130_fd_sc_hd__or3b_1 c244 (.A(net57),
    .B(net694),
    .C_N(net789),
    .X(net172));
 sky130_fd_sc_hd__nand3_2 c245 (.A(net55),
    .B(net925),
    .C(net790),
    .Y(net173));
 sky130_fd_sc_hd__and3_1 c246 (.A(net56),
    .B(net31),
    .C(net57),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 c247 (.A(net740),
    .X(net175));
 sky130_fd_sc_hd__o2111a_2 c248 (.A1(net170),
    .A2(clknet_1_0__leaf_net894),
    .B1(net925),
    .C1(net175),
    .D1(net790),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net46),
    .A1(net174),
    .A2(clknet_1_0__leaf_net921),
    .A3(net970),
    .S0(net908),
    .S1(net789),
    .X(net177));
 sky130_fd_sc_hd__and3_4 c250 (.A(net155),
    .B(net49),
    .C(clknet_1_0__leaf_net901),
    .X(net178));
 sky130_fd_sc_hd__a2111oi_1 c251 (.A1(net105),
    .A2(net178),
    .B1(net45),
    .C1(net159),
    .D1(net790),
    .Y(net179));
 sky130_fd_sc_hd__and3_1 c252 (.A(net871),
    .B(net159),
    .C(net693),
    .X(net180));
 sky130_fd_sc_hd__o2111a_4 c253 (.A1(net38),
    .A2(net173),
    .B1(net180),
    .C1(clknet_1_0__leaf_net901),
    .D1(net789),
    .X(net181));
 sky130_fd_sc_hd__or3b_2 c254 (.A(net166),
    .B(clknet_1_0__leaf_net179),
    .C_N(net958),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 c255 (.A(net740),
    .X(net183));
 sky130_fd_sc_hd__nor3b_1 c256 (.A(net183),
    .B(net175),
    .C_N(net128),
    .Y(net184));
 sky130_fd_sc_hd__mux4_4 c257 (.A0(net172),
    .A1(clknet_1_0__leaf_net179),
    .A2(net158),
    .A3(net175),
    .S0(net34),
    .S1(net790),
    .X(net185));
 sky130_fd_sc_hd__or3_1 c258 (.A(net180),
    .B(net175),
    .C(net38),
    .X(net186));
 sky130_fd_sc_hd__a2111o_1 c259 (.A1(net35),
    .A2(net186),
    .B1(net180),
    .C1(net175),
    .D1(net174),
    .X(net187));
 sky130_fd_sc_hd__inv_4 c260 (.A(net734),
    .Y(net188));
 sky130_fd_sc_hd__or3_2 c261 (.A(net175),
    .B(net188),
    .C(clknet_1_0__leaf_net776),
    .X(net920));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net128),
    .A1(net188),
    .A2(clknet_1_1__leaf_net182),
    .A3(net908),
    .S0(net919),
    .S1(clknet_1_0__leaf_net901),
    .X(net189));
 sky130_fd_sc_hd__mux4_4 c263 (.A0(net188),
    .A1(clknet_1_0__leaf_net920),
    .A2(clknet_1_0__leaf_net182),
    .A3(net970),
    .S0(net891),
    .S1(net758),
    .X(net190));
 sky130_fd_sc_hd__nand2_8 c264 (.A(net78),
    .B(net74),
    .Y(net191));
 sky130_fd_sc_hd__and2b_2 c265 (.A_N(net858),
    .B(net63),
    .X(net192));
 sky130_fd_sc_hd__nand2b_2 c266 (.A_N(net826),
    .B(net192),
    .Y(net193));
 sky130_fd_sc_hd__nor2_4 c267 (.A(net70),
    .B(net826),
    .Y(net194));
 sky130_fd_sc_hd__nand2b_1 c268 (.A_N(net76),
    .B(net194),
    .Y(net195));
 sky130_fd_sc_hd__nand2_1 c269 (.A(net831),
    .B(net66),
    .Y(net196));
 sky130_fd_sc_hd__and2b_1 c270 (.A_N(net836),
    .B(net194),
    .X(net197));
 sky130_fd_sc_hd__or2b_1 c271 (.A(net66),
    .B_N(net78),
    .X(net198));
 sky130_fd_sc_hd__nand2_2 c272 (.A(net198),
    .B(net197),
    .Y(net199));
 sky130_fd_sc_hd__nor2_2 c273 (.A(net71),
    .B(net194),
    .Y(net200));
 sky130_fd_sc_hd__or2_4 c274 (.A(net200),
    .B(net193),
    .X(net201));
 sky130_fd_sc_hd__nand3_1 c275 (.A(net191),
    .B(net71),
    .C(net201),
    .Y(net202));
 sky130_fd_sc_hd__nor3_1 c276 (.A(net197),
    .B(net74),
    .C(net869),
    .Y(net203));
 sky130_fd_sc_hd__and2_4 c277 (.A(net201),
    .B(net900),
    .X(net204));
 sky130_fd_sc_hd__or2_1 c278 (.A(net202),
    .B(net192),
    .X(net205));
 sky130_fd_sc_hd__and3_1 c279 (.A(net205),
    .B(net202),
    .C(net201),
    .X(net206));
 sky130_fd_sc_hd__nand2_1 c280 (.A(net196),
    .B(net198),
    .Y(net207));
 sky130_fd_sc_hd__or2b_1 c281 (.A(net207),
    .B_N(net205),
    .X(net208));
 sky130_fd_sc_hd__nand3_4 c282 (.A(net206),
    .B(net194),
    .C(net192),
    .Y(net896));
 sky130_fd_sc_hd__and3_1 c283 (.A(net207),
    .B(net196),
    .C(net192),
    .X(net209));
 sky130_fd_sc_hd__or2_2 c284 (.A(net193),
    .B(net209),
    .X(net210));
 sky130_fd_sc_hd__nor3b_1 c285 (.A(net195),
    .B(net208),
    .C_N(net207),
    .Y(net211));
 sky130_fd_sc_hd__nor3_1 c286 (.A(net208),
    .B(net67),
    .C(net195),
    .Y(net212));
 sky130_fd_sc_hd__and2_1 c287 (.A(net859),
    .B(net69),
    .X(net213));
 sky130_fd_sc_hd__nor2b_1 c288 (.A(net846),
    .B_N(net213),
    .Y(net214));
 sky130_fd_sc_hd__or2b_1 c289 (.A(net213),
    .B_N(net1028),
    .X(net215));
 sky130_fd_sc_hd__or4bb_4 c290 (.A(net212),
    .B(net840),
    .C_N(net79),
    .D_N(net1030),
    .X(net216));
 sky130_fd_sc_hd__nor2b_1 c291 (.A(net67),
    .B_N(net208),
    .Y(net217));
 sky130_fd_sc_hd__nand2_1 c292 (.A(net213),
    .B(net946),
    .Y(net218));
 sky130_fd_sc_hd__nor3b_1 c293 (.A(net211),
    .B(net83),
    .C_N(net831),
    .Y(net219));
 sky130_fd_sc_hd__or4bb_1 c294 (.A(net83),
    .B(net900),
    .C_N(net216),
    .D_N(net946),
    .X(net220));
 sky130_fd_sc_hd__and2b_1 c295 (.A_N(net215),
    .B(net723),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 c296 (.A(net723),
    .X(net222));
 sky130_fd_sc_hd__buf_6 c297 (.A(net723),
    .X(net223));
 sky130_fd_sc_hd__or2_1 c298 (.A(net221),
    .B(net67),
    .X(net224));
 sky130_fd_sc_hd__and3_1 c299 (.A(net65),
    .B(net223),
    .C(net722),
    .X(net225));
 sky130_fd_sc_hd__or3b_4 c300 (.A(net99),
    .B(net222),
    .C_N(net224),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__and2b_4 c302 (.A_N(net997),
    .B(net689),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 c303 (.A(net723),
    .X(net229));
 sky130_fd_sc_hd__mux4_4 c304 (.A0(net228),
    .A1(net996),
    .A2(net195),
    .A3(net225),
    .S0(net436),
    .S1(net951),
    .X(net230));
 sky130_fd_sc_hd__or3b_2 c305 (.A(net224),
    .B(net223),
    .C_N(net222),
    .X(net231));
 sky130_fd_sc_hd__sdfrtp_4 c306 (.CLK(clknet_4_0_0_clk),
    .D(net225),
    .RESET_B(net229),
    .SCD(net231),
    .SCE(net216),
    .Q(net232));
 sky130_fd_sc_hd__nor3b_1 c307 (.A(net101),
    .B(net229),
    .C_N(net231),
    .Y(net233));
 sky130_fd_sc_hd__buf_1 c308 (.A(net735),
    .X(net234));
 sky130_fd_sc_hd__nor3b_4 c309 (.A(net108),
    .B(net836),
    .C_N(net204),
    .Y(net235));
 sky130_fd_sc_hd__or3b_2 c310 (.A(net836),
    .B(net945),
    .C_N(net948),
    .X(net236));
 sky130_fd_sc_hd__and3b_1 c311 (.A_N(net852),
    .B(net222),
    .C(net120),
    .X(net237));
 sky130_fd_sc_hd__or3_4 c312 (.A(net111),
    .B(net1029),
    .C(net215),
    .X(net238));
 sky130_fd_sc_hd__o2111a_1 c313 (.A1(net870),
    .A2(net876),
    .B1(net946),
    .C1(net969),
    .D1(net722),
    .X(net239));
 sky130_fd_sc_hd__inv_2 c314 (.A(net1022),
    .Y(net240));
 sky130_fd_sc_hd__buf_16 c315 (.A(net762),
    .X(net241));
 sky130_fd_sc_hd__nor3b_4 c316 (.A(net234),
    .B(net969),
    .C_N(net743),
    .Y(net242));
 sky130_fd_sc_hd__and3_2 c317 (.A(net82),
    .B(net945),
    .C(net743),
    .X(net243));
 sky130_fd_sc_hd__inv_6 c318 (.A(net743),
    .Y(net244));
 sky130_fd_sc_hd__a2111oi_1 c319 (.A1(net222),
    .A2(net116),
    .B1(net239),
    .C1(net108),
    .D1(net788),
    .Y(net245));
 sky130_fd_sc_hd__o2111ai_1 c320 (.A1(net240),
    .A2(net242),
    .B1(net239),
    .C1(net84),
    .D1(net951),
    .Y(net246));
 sky130_fd_sc_hd__and3_1 c321 (.A(net241),
    .B(net876),
    .C(net732),
    .X(net247));
 sky130_fd_sc_hd__nor3b_2 c322 (.A(net833),
    .B(net846),
    .C_N(net222),
    .Y(net248));
 sky130_fd_sc_hd__nand3b_1 c323 (.A_N(net876),
    .B(net242),
    .C(net232),
    .Y(net249));
 sky130_fd_sc_hd__o2111a_1 c324 (.A1(net215),
    .A2(net239),
    .B1(net946),
    .C1(net945),
    .D1(net722),
    .X(net250));
 sky130_fd_sc_hd__sdfbbn_2 c325 (.CLK_N(clknet_4_2_0_clk),
    .D(net244),
    .RESET_B(net239),
    .SCD(net964),
    .SCE(net241),
    .SET_B(net743),
    .Q(net252),
    .Q_N(net251));
 sky130_fd_sc_hd__buf_2 c326 (.A(net746),
    .X(net899));
 sky130_fd_sc_hd__a2111o_4 c327 (.A1(net243),
    .A2(net238),
    .B1(clknet_1_0__leaf_net899),
    .C1(net964),
    .D1(net210),
    .X(net253));
 sky130_fd_sc_hd__a2111o_1 c328 (.A1(net945),
    .A2(net252),
    .B1(clknet_1_0__leaf_net899),
    .C1(net733),
    .D1(net763),
    .X(net254));
 sky130_fd_sc_hd__mux4_4 c329 (.A0(net230),
    .A1(net249),
    .A2(clknet_1_0__leaf_net254),
    .A3(net116),
    .S0(net862),
    .S1(net242),
    .X(net255));
 sky130_fd_sc_hd__nand2_1 c330 (.A(net232),
    .B(net252),
    .Y(net256));
 sky130_fd_sc_hd__nand2b_1 c331 (.A_N(net732),
    .B(net787),
    .Y(net257));
 sky130_fd_sc_hd__nor2_1 c332 (.A(net257),
    .B(net84),
    .Y(net258));
 sky130_fd_sc_hd__nor2b_4 c333 (.A(net106),
    .B_N(net248),
    .Y(net259));
 sky130_fd_sc_hd__and2b_1 c334 (.A_N(net134),
    .B(net734),
    .X(net260));
 sky130_fd_sc_hd__nor2_2 c335 (.A(net134),
    .B(net788),
    .Y(net261));
 sky130_fd_sc_hd__nand3b_2 c336 (.A_N(net109),
    .B(net133),
    .C(net259),
    .Y(net262));
 sky130_fd_sc_hd__or2_1 c337 (.A(net260),
    .B(net106),
    .X(net263));
 sky130_fd_sc_hd__or3_2 c338 (.A(net960),
    .B(net261),
    .C(net256),
    .X(net264));
 sky130_fd_sc_hd__nor2_1 c339 (.A(net133),
    .B(net264),
    .Y(net265));
 sky130_fd_sc_hd__or4bb_4 c340 (.A(clknet_1_0__leaf_net146),
    .B(net260),
    .C_N(net262),
    .D_N(net969),
    .X(net266));
 sky130_fd_sc_hd__or4bb_1 c341 (.A(net265),
    .B(net259),
    .C_N(net960),
    .D_N(net763),
    .X(net267));
 sky130_fd_sc_hd__or4bb_2 c342 (.A(net84),
    .B(net267),
    .C_N(net263),
    .D_N(net261),
    .X(net268));
 sky130_fd_sc_hd__sdfrtp_2 c343 (.CLK(clknet_4_9_0_clk),
    .D(net248),
    .RESET_B(net133),
    .SCD(net262),
    .SCE(net268),
    .Q(net269));
 sky130_fd_sc_hd__sdfbbn_1 c344 (.CLK_N(clknet_4_9_0_clk),
    .D(net268),
    .RESET_B(net232),
    .SCD(net248),
    .SCE(net83),
    .SET_B(net262),
    .Q(net271),
    .Q_N(net270));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net134),
    .A1(net267),
    .A2(net242),
    .A3(clknet_1_0__leaf_net143),
    .S0(net270),
    .S1(net264),
    .X(net939));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net960),
    .A1(net271),
    .A2(net900),
    .A3(net264),
    .S0(clknet_1_0__leaf_net939),
    .S1(clknet_1_0__leaf_net747),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net264),
    .A1(net271),
    .A2(net269),
    .A3(net964),
    .S0(clknet_1_0__leaf_net939),
    .S1(net259),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net265),
    .A1(net264),
    .A2(net270),
    .A3(net268),
    .S0(clknet_1_0__leaf_net939),
    .S1(net791),
    .X(net274));
 sky130_fd_sc_hd__mux4_2 c349 (.A0(net268),
    .A1(net106),
    .A2(net120),
    .A3(net270),
    .S0(clknet_1_0__leaf_net777),
    .S1(net791),
    .X(net275));
 sky130_fd_sc_hd__o2111a_2 c350 (.A1(net256),
    .A2(net960),
    .B1(net862),
    .C1(net269),
    .D1(clknet_1_0__leaf_net777),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net138),
    .A1(clknet_1_1__leaf_net146),
    .A2(net102),
    .A3(net269),
    .S0(net106),
    .S1(clknet_1_0__leaf_net777),
    .X(net277));
 sky130_fd_sc_hd__inv_1 c352 (.A(net750),
    .Y(net278));
 sky130_fd_sc_hd__and3_2 c353 (.A(clknet_1_0__leaf_net276),
    .B(net850),
    .C(net869),
    .X(net279));
 sky130_fd_sc_hd__or4bb_1 c354 (.A(net271),
    .B(net278),
    .C_N(net950),
    .D_N(net960),
    .X(net915));
 sky130_fd_sc_hd__nand3b_1 c355 (.A_N(net262),
    .B(net15),
    .C(net741),
    .Y(net280));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net120),
    .A1(net870),
    .A2(net102),
    .A3(net262),
    .S0(net280),
    .S1(net960),
    .X(net281));
 sky130_fd_sc_hd__o2111ai_2 c357 (.A1(net43),
    .A2(net878),
    .B1(net37),
    .C1(clknet_1_1__leaf_net894),
    .D1(net242),
    .Y(net933));
 sky130_fd_sc_hd__mux4_4 c358 (.A0(net258),
    .A1(net280),
    .A2(net262),
    .A3(net2),
    .S0(clknet_1_0__leaf_net153),
    .S1(clknet_1_1__leaf_net933),
    .X(net282));
 sky130_fd_sc_hd__nand3b_1 c359 (.A_N(net154),
    .B(net138),
    .C(net120),
    .Y(net928));
 sky130_fd_sc_hd__inv_2 c360 (.A(net750),
    .Y(net283));
 sky130_fd_sc_hd__or4bb_1 c361 (.A(net283),
    .B(net873),
    .C_N(net960),
    .D_N(net833),
    .X(net284));
 sky130_fd_sc_hd__mux4_2 c362 (.A0(net877),
    .A1(net138),
    .A2(net69),
    .A3(clknet_1_1__leaf_net921),
    .S0(clknet_1_1__leaf_net933),
    .S1(clknet_1_0__leaf_net939),
    .X(net285));
 sky130_fd_sc_hd__or4bb_2 c363 (.A(net138),
    .B(net271),
    .C_N(clknet_1_0__leaf_net933),
    .D_N(net43),
    .X(net286));
 sky130_fd_sc_hd__mux4_2 c364 (.A0(net149),
    .A1(clknet_1_0__leaf_net286),
    .A2(clknet_1_1__leaf_net276),
    .A3(clknet_1_0__leaf_net933),
    .S0(net43),
    .S1(clknet_1_0__leaf_net777),
    .X(net287));
 sky130_fd_sc_hd__or3b_1 c365 (.A(net37),
    .B(net960),
    .C_N(net928),
    .X(net288));
 sky130_fd_sc_hd__or4bb_4 c366 (.A(net932),
    .B(net960),
    .C_N(net30),
    .D_N(clknet_1_1__leaf_net777),
    .X(net289));
 sky130_fd_sc_hd__nand3b_4 c367 (.A_N(net867),
    .B(net154),
    .C(clknet_1_0__leaf_net289),
    .Y(net290));
 sky130_fd_sc_hd__o2111a_4 c368 (.A1(clknet_1_1__leaf_net290),
    .A2(net835),
    .B1(net138),
    .C1(net931),
    .D1(net728),
    .X(net291));
 sky130_fd_sc_hd__o2111a_2 c369 (.A1(net284),
    .A2(clknet_1_1__leaf_net290),
    .B1(clknet_1_0__leaf_net291),
    .C1(clknet_1_0__leaf_net933),
    .D1(net902),
    .X(net292));
 sky130_fd_sc_hd__mux4_4 c370 (.A0(net278),
    .A1(clknet_1_0__leaf_net290),
    .A2(net154),
    .A3(net37),
    .S0(clknet_1_0__leaf_net933),
    .S1(clknet_1_0__leaf_net291),
    .X(net293));
 sky130_fd_sc_hd__mux4_4 c371 (.A0(clknet_1_1__leaf_net153),
    .A1(clknet_1_0__leaf_net291),
    .A2(net154),
    .A3(clknet_1_0__leaf_net289),
    .S0(clknet_1_1__leaf_net292),
    .X(net294));
 sky130_fd_sc_hd__o2111a_1 c372 (.A1(net293),
    .A2(clknet_1_0__leaf_net291),
    .B1(clknet_1_1__leaf_net289),
    .C1(clknet_1_0__leaf_net290),
    .D1(clknet_1_0__leaf_net899),
    .X(net295));
 sky130_fd_sc_hd__mux4_2 c373 (.A0(net102),
    .A1(clknet_1_0__leaf_net290),
    .A2(clknet_1_0__leaf_net292),
    .A3(net900),
    .S0(net950),
    .S1(net902),
    .X(net296));
 sky130_fd_sc_hd__o2111a_1 c374 (.A1(net970),
    .A2(net932),
    .B1(net42),
    .C1(net47),
    .D1(net693),
    .X(net297));
 sky130_fd_sc_hd__o2111ai_4 c375 (.A1(clknet_1_0__leaf_net182),
    .A2(clknet_1_0__leaf_net894),
    .B1(net970),
    .C1(net694),
    .D1(clknet_1_0__leaf_net776),
    .Y(net298));
 sky130_fd_sc_hd__sdfbbp_1 c376 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_1__leaf_net291),
    .RESET_B(net173),
    .SCD(clknet_1_1__leaf_net933),
    .SCE(net47),
    .SET_B(clknet_1_1__leaf_net894),
    .Q(net300),
    .Q_N(net299));
 sky130_fd_sc_hd__or4bb_1 c377 (.A(clknet_1_1__leaf_net160),
    .B(net297),
    .C_N(net300),
    .D_N(clknet_1_1__leaf_net921),
    .X(net301));
 sky130_fd_sc_hd__nor3_4 c378 (.A(net288),
    .B(clknet_1_0__leaf_net894),
    .C(net931),
    .Y(net302));
 sky130_fd_sc_hd__a2111oi_4 c379 (.A1(net42),
    .A2(net862),
    .B1(clknet_1_0__leaf_net939),
    .C1(net844),
    .D1(clknet_1_0__leaf_net776),
    .Y(net303));
 sky130_fd_sc_hd__o2111a_1 c380 (.A1(clknet_1_1__leaf_net179),
    .A2(clknet_1_0__leaf_net302),
    .B1(clknet_1_1__leaf_net933),
    .C1(net297),
    .D1(clknet_1_0__leaf_net939),
    .X(net304));
 sky130_fd_sc_hd__o2111a_1 c381 (.A1(net188),
    .A2(clknet_1_0__leaf_net933),
    .B1(clknet_1_0__leaf_net291),
    .C1(net923),
    .D1(net728),
    .X(net924));
 sky130_fd_sc_hd__a2111oi_2 c382 (.A1(net844),
    .A2(net299),
    .B1(net875),
    .C1(clknet_1_0__leaf_net182),
    .D1(net749),
    .Y(net305));
 sky130_fd_sc_hd__or4bb_1 c383 (.A(net47),
    .B(net925),
    .C_N(clknet_1_0__leaf_net920),
    .D_N(net835),
    .X(net306));
 sky130_fd_sc_hd__mux4_2 c384 (.A0(net826),
    .A1(clknet_1_1__leaf_net302),
    .A2(net297),
    .A3(clknet_1_0__leaf_net939),
    .S0(net45),
    .S1(net299),
    .X(net307));
 sky130_fd_sc_hd__sdfbbn_2 c385 (.CLK_N(clknet_4_11_0_clk),
    .D(net300),
    .RESET_B(net908),
    .SCD(clknet_1_0__leaf_net939),
    .SCE(clknet_1_1__leaf_net747),
    .SET_B(clknet_1_1__leaf_net777),
    .Q(net309),
    .Q_N(net308));
 sky130_fd_sc_hd__mux4_4 c386 (.A0(clknet_1_1__leaf_net306),
    .A1(net948),
    .A2(clknet_1_1__leaf_net921),
    .A3(clknet_1_1__leaf_net899),
    .S0(net308),
    .S1(net733),
    .X(net310));
 sky130_fd_sc_hd__a2111oi_4 c387 (.A1(net309),
    .A2(clknet_1_1__leaf_net182),
    .B1(net128),
    .C1(clknet_1_1__leaf_net777),
    .D1(net793),
    .Y(net311));
 sky130_fd_sc_hd__mux4_4 c388 (.A0(net45),
    .A1(net42),
    .A2(net309),
    .A3(clknet_1_0__leaf_net939),
    .S0(clknet_1_0__leaf_net901),
    .S1(net793),
    .X(net312));
 sky130_fd_sc_hd__a2111o_4 c389 (.A1(net309),
    .A2(clknet_1_0__leaf_net933),
    .B1(clknet_1_1__leaf_net160),
    .C1(net878),
    .D1(net793),
    .X(net313));
 sky130_fd_sc_hd__o2111a_4 c390 (.A1(net925),
    .A2(clknet_1_1__leaf_net899),
    .B1(net774),
    .C1(clknet_1_1__leaf_net776),
    .D1(net793),
    .X(net910));
 sky130_fd_sc_hd__mux4_2 c391 (.A0(clknet_1_0__leaf_net910),
    .A1(net308),
    .A2(net740),
    .A3(net919),
    .S0(net754),
    .S1(net793),
    .X(net314));
 sky130_fd_sc_hd__mux4_4 c392 (.A0(net150),
    .A1(clknet_1_0__leaf_net306),
    .A2(net309),
    .A3(clknet_1_1__leaf_net291),
    .S0(net749),
    .S1(net793),
    .X(net315));
 sky130_fd_sc_hd__mux4_4 c393 (.A0(net55),
    .A1(clknet_1_1__leaf_net306),
    .A2(net308),
    .A3(clknet_1_1__leaf_net182),
    .S0(net889),
    .S1(net793),
    .X(net316));
 sky130_fd_sc_hd__mux4_4 c394 (.A0(net970),
    .A1(clknet_1_0__leaf_net306),
    .A2(clknet_1_0__leaf_net939),
    .A3(net740),
    .S0(net753),
    .S1(net793),
    .X(net317));
 sky130_fd_sc_hd__mux4_2 c395 (.A0(clknet_1_0__leaf_net910),
    .A1(net297),
    .A2(net753),
    .A3(net754),
    .S0(net758),
    .S1(net793),
    .X(net318));
 sky130_fd_sc_hd__nand2b_2 c396 (.A_N(net203),
    .B(net948),
    .Y(net319));
 sky130_fd_sc_hd__or2_1 c397 (.A(net338),
    .B(net900),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 c398 (.A(net686),
    .X(net321));
 sky130_fd_sc_hd__or2b_2 c399 (.A(net198),
    .B_N(net338),
    .X(net322));
 sky130_fd_sc_hd__or4bb_1 c400 (.A(net320),
    .B(net321),
    .C_N(net75),
    .D_N(net950),
    .X(net323));
 sky130_fd_sc_hd__or2_2 c401 (.A(net321),
    .B(net199),
    .X(net324));
 sky130_fd_sc_hd__and2_1 c402 (.A(net324),
    .B(net341),
    .X(net325));
 sky130_fd_sc_hd__sdfsbp_2 c403 (.CLK(clknet_4_1_0_clk),
    .D(net340),
    .SCD(net199),
    .SCE(net325),
    .SET_B(net341),
    .Q(net327),
    .Q_N(net326));
 sky130_fd_sc_hd__sdfsbp_2 c404 (.CLK(clknet_4_1_0_clk),
    .D(net206),
    .SCD(net339),
    .SCE(net326),
    .SET_B(net322),
    .Q(net329),
    .Q_N(net328));
 sky130_fd_sc_hd__inv_1 c405 (.A(net686),
    .Y(net330));
 sky130_fd_sc_hd__nor2b_2 c406 (.A(net65),
    .B_N(net199),
    .Y(net331));
 sky130_fd_sc_hd__or4bb_1 c407 (.A(net325),
    .B(net329),
    .C_N(net330),
    .D_N(net331),
    .X(net332));
 sky130_fd_sc_hd__or4bb_1 c408 (.A(net332),
    .B(net320),
    .C_N(net203),
    .D_N(net829),
    .X(net333));
 sky130_fd_sc_hd__nor3_4 c409 (.A(net324),
    .B(net326),
    .C(net686),
    .Y(net334));
 sky130_fd_sc_hd__mux4_1 c410 (.A0(net209),
    .A1(net334),
    .A2(net321),
    .A3(net79),
    .S0(net686),
    .S1(net752),
    .X(net335));
 sky130_fd_sc_hd__a2111o_1 c411 (.A1(net335),
    .A2(net898),
    .B1(net332),
    .C1(net322),
    .D1(net1019),
    .X(net336));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net331),
    .A1(net200),
    .A2(net335),
    .A3(net338),
    .S0(net752),
    .S1(net771),
    .X(net337));
 sky130_fd_sc_hd__nand2_8 c413 (.A(net193),
    .B(net131),
    .Y(net898));
 sky130_fd_sc_hd__and2_1 c414 (.A(net202),
    .B(net206),
    .X(net338));
 sky130_fd_sc_hd__and2b_4 c415 (.A_N(net77),
    .B(net885),
    .X(net339));
 sky130_fd_sc_hd__and2b_1 c416 (.A_N(net898),
    .B(net338),
    .X(net340));
 sky130_fd_sc_hd__and2_2 c417 (.A(net339),
    .B(net205),
    .X(net341));
 sky130_fd_sc_hd__nand2_2 c418 (.A(net79),
    .B(net885),
    .Y(net342));
 sky130_fd_sc_hd__inv_8 c419 (.A(net1000),
    .Y(net343));
 sky130_fd_sc_hd__clkinv_8 c420 (.A(net717),
    .Y(net344));
 sky130_fd_sc_hd__clkbuf_2 c421 (.A(net773),
    .X(net345));
 sky130_fd_sc_hd__or2b_4 c422 (.A(net72),
    .B_N(net851),
    .X(net346));
 sky130_fd_sc_hd__or3_4 c423 (.A(net343),
    .B(net65),
    .C(net967),
    .X(net347));
 sky130_fd_sc_hd__or3_1 c424 (.A(net97),
    .B(net835),
    .C(net1009),
    .X(net348));
 sky130_fd_sc_hd__mux4_2 c425 (.A0(net195),
    .A1(net226),
    .A2(net347),
    .A3(net946),
    .S0(net967),
    .S1(net689),
    .X(net349));
 sky130_fd_sc_hd__buf_16 c426 (.A(net717),
    .X(net350));
 sky130_fd_sc_hd__nand3b_1 c427 (.A_N(net838),
    .B(net201),
    .C(net967),
    .Y(net351));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(net340),
    .A1(net349),
    .A2(net966),
    .A3(net331),
    .S0(net967),
    .S1(net689),
    .X(net352));
 sky130_fd_sc_hd__sdfbbn_1 c429 (.CLK_N(clknet_4_0_0_clk),
    .D(net344),
    .RESET_B(net231),
    .SCD(net349),
    .SCE(net967),
    .SET_B(net90),
    .Q(net354),
    .Q_N(net353));
 sky130_fd_sc_hd__nand2_1 c430 (.A(net348),
    .B(net353),
    .Y(net355));
 sky130_fd_sc_hd__or3_1 c431 (.A(net229),
    .B(net354),
    .C(net966),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 c432 (.A(net717),
    .X(net357));
 sky130_fd_sc_hd__and3b_2 c433 (.A_N(net357),
    .B(net356),
    .C(net346),
    .X(net358));
 sky130_fd_sc_hd__and3b_1 c434 (.A_N(net354),
    .B(net191),
    .C(net358),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net359),
    .A1(net85),
    .A2(net950),
    .A3(net90),
    .S0(net349),
    .S1(net353),
    .X(net360));
 sky130_fd_sc_hd__a2111oi_1 c436 (.A1(net355),
    .A2(net356),
    .B1(net358),
    .C1(net967),
    .D1(net966),
    .Y(net361));
 sky130_fd_sc_hd__o2111ai_1 c437 (.A1(net356),
    .A2(net213),
    .B1(net340),
    .C1(net967),
    .D1(net946),
    .Y(net362));
 sky130_fd_sc_hd__o2111a_4 c438 (.A1(net359),
    .A2(net343),
    .B1(net97),
    .C1(net721),
    .D1(clknet_1_0__leaf_net794),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net967),
    .A1(net361),
    .A2(net97),
    .A3(net835),
    .S0(net359),
    .S1(net721),
    .X(net364));
 sky130_fd_sc_hd__or3b_2 c440 (.A(net237),
    .B(net251),
    .C_N(clknet_1_0__leaf_net794),
    .X(net365));
 sky130_fd_sc_hd__a2111o_2 c441 (.A1(net75),
    .A2(clknet_1_0__leaf_net365),
    .B1(net950),
    .C1(clknet_1_0__leaf_net899),
    .D1(net689),
    .X(net366));
 sky130_fd_sc_hd__buf_6 c442 (.A(net681),
    .X(net367));
 sky130_fd_sc_hd__a2111o_4 c443 (.A1(net851),
    .A2(net72),
    .B1(clknet_1_0__leaf_net899),
    .C1(net122),
    .D1(net97),
    .X(net368));
 sky130_fd_sc_hd__o2111ai_4 c444 (.A1(net126),
    .A2(net898),
    .B1(net347),
    .C1(net946),
    .D1(clknet_1_0__leaf_net794),
    .Y(net369));
 sky130_fd_sc_hd__nand3_2 c445 (.A(net364),
    .B(net2),
    .C(net946),
    .Y(net370));
 sky130_fd_sc_hd__nor3b_1 c446 (.A(clknet_1_0__leaf_net365),
    .B(net341),
    .C_N(net947),
    .Y(net371));
 sky130_fd_sc_hd__or3_4 c447 (.A(net368),
    .B(net346),
    .C(net951),
    .X(net372));
 sky130_fd_sc_hd__and3b_1 c448 (.A_N(net878),
    .B(clknet_1_0__leaf_net372),
    .C(net689),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net349),
    .A1(net948),
    .A2(net953),
    .A3(net945),
    .S0(net342),
    .S1(net951),
    .X(net374));
 sky130_fd_sc_hd__nor2b_1 c450 (.A(net232),
    .B_N(net75),
    .Y(net375));
 sky130_fd_sc_hd__inv_4 c451 (.A(net681),
    .Y(net376));
 sky130_fd_sc_hd__buf_6 c452 (.A(net717),
    .X(net907));
 sky130_fd_sc_hd__inv_1 c453 (.A(net723),
    .Y(net377));
 sky130_fd_sc_hd__or4bb_2 c454 (.A(net341),
    .B(net339),
    .C_N(net346),
    .D_N(net377),
    .X(net378));
 sky130_fd_sc_hd__nor2b_1 c455 (.A(clknet_1_0__leaf_net372),
    .B_N(net378),
    .Y(net379));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net85),
    .A1(net875),
    .A2(clknet_1_0__leaf_net379),
    .A3(clknet_1_0__leaf_net365),
    .S0(net342),
    .S1(net771),
    .X(net380));
 sky130_fd_sc_hd__mux4_2 c457 (.A0(net377),
    .A1(net232),
    .A2(net343),
    .A3(net341),
    .S0(net375),
    .S1(net682),
    .X(net381));
 sky130_fd_sc_hd__a2111o_4 c458 (.A1(net946),
    .A2(clknet_1_0__leaf_net366),
    .B1(net850),
    .C1(net381),
    .D1(net682),
    .X(net382));
 sky130_fd_sc_hd__sdfbbp_1 c459 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_1__leaf_net379),
    .RESET_B(net238),
    .SCD(net370),
    .SCE(net376),
    .SET_B(net1010),
    .Q(net886),
    .Q_N(net383));
 sky130_fd_sc_hd__mux4_2 c460 (.A0(net370),
    .A1(net334),
    .A2(net381),
    .A3(clknet_1_0__leaf_net373),
    .S0(clknet_1_0__leaf_net366),
    .S1(net1025),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net381),
    .A1(net236),
    .A2(net886),
    .A3(net1020),
    .S0(net771),
    .S1(net1016),
    .X(net385));
 sky130_fd_sc_hd__nand3b_4 c462 (.A_N(net263),
    .B(net347),
    .C(net1026),
    .Y(net386));
 sky130_fd_sc_hd__or4bb_1 c463 (.A(net948),
    .B(net763),
    .C_N(net791),
    .D_N(clknet_1_0__leaf_net794),
    .X(net387));
 sky130_fd_sc_hd__buf_4 c464 (.A(net735),
    .X(net930));
 sky130_fd_sc_hd__or4bb_1 c465 (.A(net375),
    .B(net1025),
    .C_N(net386),
    .D_N(net1010),
    .X(net388));
 sky130_fd_sc_hd__or4bb_4 c466 (.A(net147),
    .B(net191),
    .C_N(clknet_1_0__leaf_net747),
    .D_N(net347),
    .X(net389));
 sky130_fd_sc_hd__or4bb_1 c467 (.A(net129),
    .B(net259),
    .C_N(net930),
    .D_N(net263),
    .X(net390));
 sky130_fd_sc_hd__or3_1 c468 (.A(net347),
    .B(net930),
    .C(net261),
    .X(net391));
 sky130_fd_sc_hd__sdfbbn_1 c469 (.CLK_N(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net387),
    .RESET_B(net269),
    .SCD(net390),
    .SCE(net388),
    .SET_B(net263),
    .Q(net393),
    .Q_N(net392));
 sky130_fd_sc_hd__mux4_2 c470 (.A0(net390),
    .A1(clknet_1_1__leaf_net389),
    .A2(net392),
    .A3(net383),
    .S0(net122),
    .S1(net911),
    .X(net394));
 sky130_fd_sc_hd__a2111o_2 c471 (.A1(clknet_1_1__leaf_net143),
    .A2(net129),
    .B1(net393),
    .C1(net930),
    .D1(net992),
    .X(net395));
 sky130_fd_sc_hd__sdfbbn_2 c472 (.CLK_N(clknet_4_12_0_clk),
    .D(net269),
    .RESET_B(net388),
    .SCD(net259),
    .SCE(net930),
    .SET_B(clknet_1_1__leaf_net939),
    .Q(net916),
    .Q_N(net396));
 sky130_fd_sc_hd__or4bb_4 c473 (.A(net367),
    .B(net391),
    .C_N(clknet_1_0__leaf_net939),
    .D_N(net191),
    .X(net397));
 sky130_fd_sc_hd__a2111o_2 c474 (.A1(net393),
    .A2(net916),
    .B1(net261),
    .C1(clknet_1_0__leaf_net394),
    .D1(clknet_1_0__leaf_net747),
    .X(net398));
 sky130_fd_sc_hd__or4bb_4 c475 (.A(clknet_1_0__leaf_net389),
    .B(net973),
    .C_N(net269),
    .D_N(net763),
    .X(net399));
 sky130_fd_sc_hd__or4bb_2 c476 (.A(clknet_1_1__leaf_net394),
    .B(net259),
    .C_N(net700),
    .D_N(net1026),
    .X(net400));
 sky130_fd_sc_hd__a2111oi_0 c477 (.A1(net388),
    .A2(net337),
    .B1(net261),
    .C1(net347),
    .D1(clknet_1_0__leaf_net373),
    .Y(net401));
 sky130_fd_sc_hd__sdfstp_2 c478 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net899),
    .SCD(clknet_1_1__leaf_net939),
    .SCE(net1023),
    .SET_B(net1013),
    .Q(net402));
 sky130_fd_sc_hd__sdfstp_1 c479 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net387),
    .SCD(net869),
    .SCE(net968),
    .SET_B(clknet_1_0__leaf_net747),
    .Q(net403));
 sky130_fd_sc_hd__or4bb_1 c480 (.A(net147),
    .B(net973),
    .C_N(net916),
    .D_N(net82),
    .X(net404));
 sky130_fd_sc_hd__mux4_2 c481 (.A0(net930),
    .A1(net232),
    .A2(net402),
    .A3(clknet_1_0__leaf_net394),
    .S0(net699),
    .S1(net780),
    .X(net405));
 sky130_fd_sc_hd__or4bb_4 c482 (.A(net404),
    .B(net991),
    .C_N(net780),
    .D_N(clknet_1_0__leaf_net795),
    .X(net406));
 sky130_fd_sc_hd__mux4_4 c483 (.A0(clknet_1_1__leaf_net406),
    .A1(net403),
    .A2(net404),
    .A3(clknet_1_0__leaf_net399),
    .S0(net973),
    .S1(net392),
    .X(net407));
 sky130_fd_sc_hd__or4bb_1 c484 (.A(net391),
    .B(net123),
    .C_N(clknet_1_1__leaf_net254),
    .D_N(net796),
    .X(net408));
 sky130_fd_sc_hd__nor3_4 c485 (.A(net422),
    .B(clknet_1_1__leaf_net289),
    .C(clknet_1_1__leaf_net748),
    .Y(net937));
 sky130_fd_sc_hd__inv_2 c486 (.A(net772),
    .Y(net409));
 sky130_fd_sc_hd__clkbuf_2 c487 (.A(net772),
    .X(net410));
 sky130_fd_sc_hd__nand3_1 c488 (.A(net378),
    .B(net422),
    .C(net896),
    .Y(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 c489 (.A(clknet_1_1__leaf_net748),
    .X(net412));
 sky130_fd_sc_hd__inv_6 c490 (.A(net735),
    .Y(net897));
 sky130_fd_sc_hd__nor3b_1 c491 (.A(net409),
    .B(net386),
    .C_N(net931),
    .Y(net929));
 sky130_fd_sc_hd__inv_4 c492 (.A(net727),
    .Y(net413));
 sky130_fd_sc_hd__nor3b_2 c493 (.A(net412),
    .B(net986),
    .C_N(net897),
    .Y(net414));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(clknet_1_1__leaf_net161),
    .A1(net411),
    .A2(net409),
    .A3(net383),
    .S0(clknet_1_1__leaf_net795),
    .S1(net796),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 c495 (.A(net727),
    .X(net416));
 sky130_fd_sc_hd__mux4_4 c496 (.A0(net416),
    .A1(clknet_1_0__leaf_net937),
    .A2(net896),
    .A3(net410),
    .S0(net898),
    .S1(clknet_1_1__leaf_net423),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net163),
    .A1(clknet_1_1__leaf_net286),
    .A2(net985),
    .A3(net416),
    .S0(net396),
    .S1(net759),
    .X(net418));
 sky130_fd_sc_hd__mux4_4 c498 (.A0(clknet_1_1__leaf_net366),
    .A1(net984),
    .A2(clknet_1_0__leaf_net414),
    .A3(net410),
    .S0(clknet_1_0__leaf_net748),
    .S1(net759),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net419),
    .A1(net422),
    .A2(clknet_1_1__leaf_net425),
    .A3(net886),
    .S0(clknet_1_0__leaf_net904),
    .S1(net935),
    .X(net420));
 sky130_fd_sc_hd__or2b_1 c500 (.A(net436),
    .B_N(net771),
    .X(net421));
 sky130_fd_sc_hd__inv_2 c201_13 (.A(clknet_1_1__leaf_net776),
    .Y(net987));
 sky130_fd_sc_hd__or4bb_4 c502 (.A(net2),
    .B(net931),
    .C_N(net421),
    .D_N(net923),
    .X(net422));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net422),
    .A1(net983),
    .A2(net261),
    .A3(net966),
    .S0(clknet_1_1__leaf_net366),
    .S1(net383),
    .X(net423));
 sky130_fd_sc_hd__mux4_2 c504 (.A0(clknet_1_0__leaf_net286),
    .A1(net842),
    .A2(net990),
    .A3(net923),
    .S0(net422),
    .S1(net982),
    .X(net424));
 sky130_fd_sc_hd__and3b_1 c505 (.A_N(net261),
    .B(clknet_1_0__leaf_net795),
    .C(net935),
    .X(net425));
 sky130_fd_sc_hd__mux4_4 c526 (.A0(net49),
    .A1(clknet_1_0__leaf_net289),
    .A2(net869),
    .A3(net927),
    .S0(net934),
    .S1(net922),
    .X(net914));
 sky130_fd_sc_hd__mux4_2 c527 (.A0(net912),
    .A1(clknet_1_0__leaf_net924),
    .A2(net966),
    .A3(net936),
    .S0(net889),
    .S1(clknet_1_1__leaf_net795),
    .X(net426));
 sky130_fd_sc_hd__or2b_1 c528 (.A(net196),
    .B_N(net331),
    .X(net427));
 sky130_fd_sc_hd__nand2_1 c529 (.A(net205),
    .B(net329),
    .Y(net428));
 sky130_fd_sc_hd__and2_1 c530 (.A(net338),
    .B(net200),
    .X(net429));
 sky130_fd_sc_hd__nor3b_1 c531 (.A(net82),
    .B(net334),
    .C_N(net771),
    .Y(net430));
 sky130_fd_sc_hd__nand2_1 c532 (.A(net325),
    .B(net330),
    .Y(net431));
 sky130_fd_sc_hd__or3b_1 c533 (.A(net325),
    .B(net943),
    .C_N(net771),
    .X(net432));
 sky130_fd_sc_hd__inv_2 c534 (.A(net685),
    .Y(net433));
 sky130_fd_sc_hd__clkbuf_8 c535 (.A(net746),
    .X(net434));
 sky130_fd_sc_hd__nand2b_1 c536 (.A_N(net427),
    .B(net943),
    .Y(net435));
 sky130_fd_sc_hd__clkinv_2 c501_4 (.A(clknet_1_1__leaf_net748),
    .Y(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 c538 (.A(net761),
    .X(net437));
 sky130_fd_sc_hd__and2_1 c539 (.A(net943),
    .B(net434),
    .X(net438));
 sky130_fd_sc_hd__or2b_4 c540 (.A(net437),
    .B_N(net977),
    .X(net439));
 sky130_fd_sc_hd__nor3b_1 c541 (.A(net330),
    .B(net976),
    .C_N(net950),
    .Y(net440));
 sky130_fd_sc_hd__buf_6 c542 (.A(net761),
    .X(net441));
 sky130_fd_sc_hd__dlymetal6s2s_1 c543 (.A(net746),
    .X(net442));
 sky130_fd_sc_hd__inv_2 c544 (.A(net685),
    .Y(net443));
 sky130_fd_sc_hd__o2111a_2 c545 (.A1(net975),
    .A2(clknet_1_1__leaf_net442),
    .B1(net941),
    .C1(net82),
    .D1(net943),
    .X(net444));
 sky130_fd_sc_hd__nor2_2 c546 (.A(net443),
    .B(clknet_1_0__leaf_net442),
    .Y(net445));
 sky130_fd_sc_hd__and2b_1 c547 (.A_N(net428),
    .B(net685),
    .X(net446));
 sky130_fd_sc_hd__nor3_2 c548 (.A(net324),
    .B(clknet_1_0__leaf_net440),
    .C(clknet_1_0__leaf_net445),
    .Y(net447));
 sky130_fd_sc_hd__inv_1 c549 (.A(net761),
    .Y(net448));
 sky130_fd_sc_hd__and3_1 c550 (.A(net90),
    .B(net344),
    .C(net946),
    .X(net449));
 sky130_fd_sc_hd__nor3b_1 c551 (.A(net344),
    .B(net948),
    .C_N(net943),
    .Y(net450));
 sky130_fd_sc_hd__nand3_4 c552 (.A(net448),
    .B(net943),
    .C(net344),
    .Y(net451));
 sky130_fd_sc_hd__or3b_1 c553 (.A(net357),
    .B(net943),
    .C_N(clknet_1_0__leaf_net363),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 c554 (.A(net765),
    .X(net453));
 sky130_fd_sc_hd__clkinv_4 c555 (.A(net765),
    .Y(net454));
 sky130_fd_sc_hd__nand3b_4 c556 (.A_N(net829),
    .B(net201),
    .C(net454),
    .Y(net455));
 sky130_fd_sc_hd__a2111o_4 c557 (.A1(clknet_1_0__leaf_net452),
    .A2(net450),
    .B1(net943),
    .C1(clknet_1_0__leaf_net363),
    .D1(clknet_1_1__leaf_net794),
    .X(net456));
 sky130_fd_sc_hd__or2b_1 c558 (.A(net331),
    .B_N(net344),
    .X(net457));
 sky130_fd_sc_hd__o2111ai_4 c559 (.A1(net449),
    .A2(clknet_1_0__leaf_net445),
    .B1(net973),
    .C1(net358),
    .D1(net451),
    .Y(net458));
 sky130_fd_sc_hd__and3b_2 c560 (.A_N(net95),
    .B(net453),
    .C(net201),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net457),
    .A1(clknet_1_0__leaf_net445),
    .A2(net459),
    .A3(net943),
    .S0(clknet_1_0__leaf_net363),
    .S1(net357),
    .X(net460));
 sky130_fd_sc_hd__o2111a_1 c562 (.A1(clknet_1_0__leaf_net460),
    .A2(net327),
    .B1(net459),
    .C1(net944),
    .D1(net1001),
    .X(net461));
 sky130_fd_sc_hd__mux4_4 c563 (.A0(clknet_1_1__leaf_net460),
    .A1(clknet_1_1__leaf_net452),
    .A2(net455),
    .A3(net459),
    .S0(net684),
    .S1(net774),
    .X(net462));
 sky130_fd_sc_hd__or3b_2 c564 (.A(net459),
    .B(net900),
    .C_N(net448),
    .X(net463));
 sky130_fd_sc_hd__nand3b_2 c565 (.A_N(net344),
    .B(net357),
    .C(net782),
    .Y(net464));
 sky130_fd_sc_hd__buf_1 c566 (.A(net720),
    .X(net465));
 sky130_fd_sc_hd__sdfbbp_1 c567 (.CLK(clknet_4_1_0_clk),
    .D(net457),
    .RESET_B(net459),
    .SCD(net455),
    .SCE(net941),
    .SET_B(net782),
    .Q(net467),
    .Q_N(net466));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net358),
    .A1(net464),
    .A2(net319),
    .A3(net944),
    .S0(net941),
    .S1(net684),
    .X(net468));
 sky130_fd_sc_hd__o2111ai_4 c569 (.A1(net465),
    .A2(net459),
    .B1(net467),
    .C1(net334),
    .D1(net463),
    .Y(net469));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net201),
    .A1(net451),
    .A2(net455),
    .A3(net1014),
    .S0(net782),
    .S1(net797),
    .X(net470));
 sky130_fd_sc_hd__mux4_4 c571 (.A0(net450),
    .A1(net950),
    .A2(net465),
    .A3(net463),
    .S0(net346),
    .S1(net466),
    .X(net471));
 sky130_fd_sc_hd__o2111a_4 c572 (.A1(net464),
    .A2(net455),
    .B1(clknet_1_0__leaf_net440),
    .C1(net453),
    .D1(net951),
    .X(net472));
 sky130_fd_sc_hd__sdfstp_2 c573 (.CLK(clknet_4_1_0_clk),
    .D(clknet_1_1__leaf_net445),
    .SCD(net337),
    .SCE(net967),
    .SET_B(net1015),
    .Q(net473));
 sky130_fd_sc_hd__o2111a_1 c574 (.A1(net337),
    .A2(net464),
    .B1(net383),
    .C1(net204),
    .D1(net798),
    .X(net474));
 sky130_fd_sc_hd__o2111ai_4 c575 (.A1(net467),
    .A2(net907),
    .B1(net952),
    .C1(net473),
    .D1(net800),
    .Y(net475));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net455),
    .A1(net454),
    .A2(net343),
    .A3(net966),
    .S0(net751),
    .S1(net887),
    .X(net476));
 sky130_fd_sc_hd__o2111ai_1 c577 (.A1(net343),
    .A2(net476),
    .B1(clknet_1_0__leaf_net440),
    .C1(net72),
    .D1(net797),
    .Y(net477));
 sky130_fd_sc_hd__or4bb_1 c578 (.A(clknet_1_1__leaf_net440),
    .B(net968),
    .C_N(net473),
    .D_N(net751),
    .X(net478));
 sky130_fd_sc_hd__sdfbbn_2 c579 (.CLK_N(clknet_4_3_0_clk),
    .D(net476),
    .RESET_B(net475),
    .SCD(clknet_1_0__leaf_net371),
    .SCE(clknet_1_1__leaf_net372),
    .SET_B(net473),
    .Q(net480),
    .Q_N(net479));
 sky130_fd_sc_hd__sdfbbn_2 c580 (.CLK_N(clknet_4_6_0_clk),
    .D(net475),
    .RESET_B(clknet_1_0__leaf_net373),
    .SCD(clknet_1_0__leaf_net477),
    .SCE(clknet_1_1__leaf_net445),
    .SET_B(net346),
    .Q(net938),
    .Q_N(net481));
 sky130_fd_sc_hd__sdfbbp_1 c581 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net371),
    .RESET_B(clknet_1_0__leaf_net366),
    .SCD(net466),
    .SCE(net251),
    .SET_B(net683),
    .Q(net483),
    .Q_N(net482));
 sky130_fd_sc_hd__a2111o_2 c582 (.A1(clknet_1_1__leaf_net478),
    .A2(net950),
    .B1(clknet_1_1__leaf_net440),
    .C1(net482),
    .D1(clknet_1_0__leaf_net382),
    .X(net484));
 sky130_fd_sc_hd__o2111ai_2 c583 (.A1(clknet_1_0__leaf_net472),
    .A2(clknet_1_0__leaf_net372),
    .B1(net337),
    .C1(net473),
    .D1(net479),
    .Y(net485));
 sky130_fd_sc_hd__or4bb_4 c584 (.A(clknet_1_1__leaf_net382),
    .B(net473),
    .C_N(net903),
    .D_N(clknet_1_1__leaf_net794),
    .X(net486));
 sky130_fd_sc_hd__a2111oi_2 c585 (.A1(net453),
    .A2(net339),
    .B1(net479),
    .C1(clknet_1_0__leaf_net472),
    .D1(net775),
    .Y(net487));
 sky130_fd_sc_hd__or4bb_1 c586 (.A(net346),
    .B(net482),
    .C_N(net756),
    .D_N(net775),
    .X(net488));
 sky130_fd_sc_hd__o2111ai_2 c587 (.A1(net488),
    .A2(net480),
    .B1(net204),
    .C1(net123),
    .D1(net467),
    .Y(net489));
 sky130_fd_sc_hd__mux4_4 c588 (.A0(clknet_1_1__leaf_net477),
    .A1(clknet_1_0__leaf_net472),
    .A2(net941),
    .A3(clknet_1_1__leaf_net373),
    .S0(net913),
    .S1(net775),
    .X(net490));
 sky130_fd_sc_hd__o2111a_4 c589 (.A1(net334),
    .A2(net475),
    .B1(net489),
    .C1(net467),
    .D1(net799),
    .X(net892));
 sky130_fd_sc_hd__mux4_2 c590 (.A0(net938),
    .A1(net473),
    .A2(net251),
    .A3(clknet_1_1__leaf_net440),
    .S0(net892),
    .S1(net756),
    .X(net491));
 sky130_fd_sc_hd__sdfbbn_2 c591 (.CLK_N(clknet_4_6_0_clk),
    .D(net238),
    .RESET_B(net892),
    .SCD(net346),
    .SCE(clknet_1_1__leaf_net372),
    .SET_B(net1018),
    .Q(net493),
    .Q_N(net492));
 sky130_fd_sc_hd__mux4_4 c592 (.A0(clknet_1_1__leaf_net372),
    .A1(net892),
    .A2(net204),
    .A3(net492),
    .S0(net903),
    .S1(net906),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net489),
    .A1(net945),
    .A2(clknet_1_0__leaf_net478),
    .A3(clknet_1_0__leaf_net472),
    .S0(net826),
    .S1(net892),
    .X(net495));
 sky130_fd_sc_hd__sedfxbp_1 c594 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net472),
    .DE(net826),
    .SCD(clknet_1_0__leaf_net517),
    .SCE(net762),
    .Q(net497),
    .Q_N(net496));
 sky130_fd_sc_hd__a2111o_1 c595 (.A1(clknet_1_1__leaf_net516),
    .A2(net941),
    .B1(clknet_1_1__leaf_net373),
    .C1(net259),
    .D1(net764),
    .X(net498));
 sky130_fd_sc_hd__o2111ai_1 c596 (.A1(net473),
    .A2(net123),
    .B1(net511),
    .C1(clknet_1_0__leaf_net517),
    .D1(net911),
    .Y(net499));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net123),
    .A1(net952),
    .A2(net945),
    .A3(net683),
    .S0(net762),
    .S1(net764),
    .X(net500));
 sky130_fd_sc_hd__mux4_2 c598 (.A0(clknet_1_1__leaf_net373),
    .A1(net488),
    .A2(clknet_1_0__leaf_net516),
    .A3(net328),
    .S0(net973),
    .S1(net754),
    .X(net501));
 sky130_fd_sc_hd__sdfbbn_1 c599 (.CLK_N(clknet_4_12_0_clk),
    .D(net941),
    .RESET_B(net514),
    .SCD(net511),
    .SCE(clknet_1_0__leaf_net407),
    .SET_B(net803),
    .Q(net503),
    .Q_N(net502));
 sky130_fd_sc_hd__or4bb_1 c600 (.A(net510),
    .B(net519),
    .C_N(net339),
    .D_N(net513),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net128),
    .A1(net504),
    .A2(net403),
    .A3(clknet_1_0__leaf_net517),
    .S0(net513),
    .S1(net803),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net500),
    .A1(net504),
    .A2(net496),
    .A3(net754),
    .S0(net786),
    .S1(net797),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net510),
    .A1(net504),
    .A2(net500),
    .A3(net496),
    .S0(net791),
    .S1(net804),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net500),
    .A1(net504),
    .A2(clknet_1_0__leaf_net407),
    .A3(net886),
    .S0(net760),
    .S1(net804),
    .X(net508));
 sky130_fd_sc_hd__a2111oi_1 c605 (.A1(net973),
    .A2(net454),
    .B1(net492),
    .C1(net403),
    .D1(net800),
    .Y(net509));
 sky130_fd_sc_hd__mux4_4 c606 (.A0(net403),
    .A1(clknet_1_0__leaf_net366),
    .A2(net93),
    .A3(net339),
    .S0(net903),
    .S1(net798),
    .X(net917));
 sky130_fd_sc_hd__a2111o_1 c607 (.A1(net375),
    .A2(net857),
    .B1(net252),
    .C1(net967),
    .D1(net840),
    .X(net510));
 sky130_fd_sc_hd__sedfxbp_1 c608 (.CLK(clknet_4_3_0_clk),
    .D(net93),
    .DE(net941),
    .SCD(net337),
    .SCE(clknet_1_0__leaf_net794),
    .Q(net512),
    .Q_N(net511));
 sky130_fd_sc_hd__sdfbbp_1 c609 (.CLK(clknet_4_3_0_clk),
    .D(net941),
    .RESET_B(net1017),
    .SCD(net386),
    .SCE(net93),
    .SET_B(net1012),
    .Q(net514),
    .Q_N(net513));
 sky130_fd_sc_hd__or4bb_1 c610 (.A(net346),
    .B(net968),
    .C_N(net513),
    .D_N(net906),
    .X(net515));
 sky130_fd_sc_hd__mux4_2 c611 (.A0(net512),
    .A1(clknet_1_0__leaf_net406),
    .A2(net396),
    .A3(net481),
    .S0(net774),
    .S1(net798),
    .X(net516));
 sky130_fd_sc_hd__or4bb_1 c612 (.A(net1005),
    .B(net454),
    .C_N(clknet_1_0__leaf_net516),
    .D_N(net799),
    .X(net517));
 sky130_fd_sc_hd__sdfbbn_2 c613 (.CLK_N(clknet_4_3_0_clk),
    .D(net963),
    .RESET_B(clknet_1_0__leaf_net517),
    .SCD(net840),
    .SCE(net455),
    .SET_B(net798),
    .Q(net519),
    .Q_N(net518));
 sky130_fd_sc_hd__a2111oi_1 c614 (.A1(net339),
    .A2(net938),
    .B1(net514),
    .C1(net429),
    .D1(net1021),
    .Y(net520));
 sky130_fd_sc_hd__mux4_2 c615 (.A0(net514),
    .A1(net402),
    .A2(clknet_1_1__leaf_net516),
    .A3(clknet_1_0__leaf_net917),
    .S0(net913),
    .S1(net802),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net123),
    .A1(net30),
    .A2(net518),
    .A3(net252),
    .S0(net502),
    .S1(net753),
    .X(net522));
 sky130_fd_sc_hd__mux4_4 c617 (.A0(net454),
    .A1(net252),
    .A2(clknet_1_0__leaf_net414),
    .A3(net163),
    .S0(net792),
    .S1(clknet_1_0__leaf_net904),
    .X(net523));
 sky130_fd_sc_hd__mux4_4 c618 (.A0(clknet_1_1__leaf_net366),
    .A1(net966),
    .A2(net163),
    .A3(net981),
    .S0(net251),
    .S1(net792),
    .X(net524));
 sky130_fd_sc_hd__mux4_4 c619 (.A0(net413),
    .A1(net892),
    .A2(net515),
    .A3(clknet_1_1__leaf_net414),
    .S0(net251),
    .S1(net792),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c62 (.A0(net828),
    .A1(net866),
    .A2(net839),
    .A3(net845),
    .S0(net867),
    .S1(net856),
    .X(net0));
 sky130_fd_sc_hd__mux4_4 c620 (.A0(net163),
    .A1(clknet_1_1__leaf_net899),
    .A2(net128),
    .A3(net913),
    .S0(net887),
    .S1(clknet_1_0__leaf_net904),
    .X(net526));
 sky130_fd_sc_hd__mux4_2 c621 (.A0(net252),
    .A1(net519),
    .A2(net958),
    .A3(clknet_1_1__leaf_net366),
    .S0(net402),
    .S1(net951),
    .X(net527));
 sky130_fd_sc_hd__mux4_2 c622 (.A0(net410),
    .A1(net844),
    .A2(net519),
    .A3(net327),
    .S0(net966),
    .S1(net907),
    .X(net888));
 sky130_fd_sc_hd__mux4_2 c623 (.A0(net30),
    .A1(net523),
    .A2(clknet_1_1__leaf_net939),
    .A3(clknet_1_0__leaf_net527),
    .S0(net413),
    .S1(net808),
    .X(net528));
 sky130_fd_sc_hd__mux4_2 c624 (.A0(net402),
    .A1(clknet_1_0__leaf_net527),
    .A2(net503),
    .A3(net989),
    .S0(net518),
    .S1(net909),
    .X(net529));
 sky130_fd_sc_hd__mux4_4 c625 (.A0(net480),
    .A1(net128),
    .A2(net31),
    .A3(net792),
    .S0(net805),
    .S1(net808),
    .X(net530));
 sky130_fd_sc_hd__mux4_4 c626 (.A0(clknet_1_1__leaf_net414),
    .A1(clknet_1_1__leaf_net527),
    .A2(net454),
    .A3(net386),
    .S0(net753),
    .S1(net760),
    .X(net531));
 sky130_fd_sc_hd__mux4_4 c627 (.A0(net163),
    .A1(net952),
    .A2(net402),
    .A3(net980),
    .S0(net700),
    .S1(net810),
    .X(net905));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net833),
    .A1(net454),
    .A2(clknet_1_1__leaf_net527),
    .A3(net888),
    .S0(net760),
    .S1(net810),
    .X(net532));
 sky130_fd_sc_hd__mux4_4 c629 (.A0(net503),
    .A1(net454),
    .A2(clknet_1_1__leaf_net527),
    .A3(net806),
    .S0(net807),
    .S1(net809),
    .X(net533));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net0),
    .A1(net862),
    .A2(net839),
    .A3(net856),
    .S0(net866),
    .S1(net867),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net402),
    .A1(net907),
    .A2(net988),
    .A3(net806),
    .S0(net809),
    .S1(net810),
    .X(net534));
 sky130_fd_sc_hd__mux4_4 c631 (.A0(net515),
    .A1(net534),
    .A2(clknet_1_1__leaf_net414),
    .A3(net805),
    .S0(net807),
    .S1(net809),
    .X(net893));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net31),
    .A1(net455),
    .A2(net850),
    .A3(net30),
    .S0(net772),
    .S1(net809),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net522),
    .A1(net502),
    .A2(net897),
    .A3(net887),
    .S0(net802),
    .S1(net810),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net163),
    .A1(net938),
    .A2(net123),
    .A3(clknet_1_1__leaf_net899),
    .S0(clknet_1_0__leaf_net527),
    .S1(net888),
    .X(net537));
 sky130_fd_sc_hd__mux4_2 c635 (.A0(net536),
    .A1(net535),
    .A2(net31),
    .A3(net122),
    .S0(clknet_1_0__leaf_net905),
    .S1(net807),
    .X(net538));
 sky130_fd_sc_hd__mux4_2 c636 (.A0(net455),
    .A1(net480),
    .A2(clknet_1_1__leaf_net527),
    .A3(net951),
    .S0(net772),
    .S1(net808),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net916),
    .A1(net979),
    .A2(net760),
    .A3(net774),
    .S0(clknet_1_0__leaf_net904),
    .S1(net810),
    .X(net540));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net839),
    .A1(net882),
    .A2(net867),
    .A3(net863),
    .S0(net878),
    .S1(net1),
    .X(net2));
 sky130_fd_sc_hd__mux4_1 c65 (.A0(net856),
    .A1(net835),
    .A2(net849),
    .A3(net826),
    .S0(net851),
    .S1(net857),
    .X(net3));
 sky130_fd_sc_hd__or2_1 c66 (.A(net0),
    .B(net879),
    .X(net4));
 sky130_fd_sc_hd__or2_1 c660 (.A(net557),
    .B(net326),
    .X(net541));
 sky130_fd_sc_hd__and2_4 c661 (.A(net561),
    .B(net199),
    .X(net542));
 sky130_fd_sc_hd__or2_2 c662 (.A(net199),
    .B(net542),
    .X(net543));
 sky130_fd_sc_hd__or2b_1 c663 (.A(net847),
    .B_N(net965),
    .X(net544));
 sky130_fd_sc_hd__or2b_1 c664 (.A(clknet_1_1__leaf_net439),
    .B_N(net194),
    .X(net545));
 sky130_fd_sc_hd__and2b_2 c665 (.A_N(net560),
    .B(net869),
    .X(net546));
 sky130_fd_sc_hd__or2b_1 c666 (.A(net557),
    .B_N(net962),
    .X(net547));
 sky130_fd_sc_hd__nand2_2 c667 (.A(net559),
    .B(net543),
    .Y(net548));
 sky130_fd_sc_hd__or2b_1 c668 (.A(net204),
    .B_N(net548),
    .X(net549));
 sky130_fd_sc_hd__nand2b_1 c669 (.A_N(net544),
    .B(net557),
    .Y(net550));
 sky130_fd_sc_hd__nor2b_1 c67 (.A(net841),
    .B_N(net863),
    .Y(net5));
 sky130_fd_sc_hd__nor3b_1 c670 (.A(net548),
    .B(clknet_1_1__leaf_net447),
    .C_N(net558),
    .Y(net551));
 sky130_fd_sc_hd__nand3b_4 c671 (.A_N(net545),
    .B(net548),
    .C(net962),
    .Y(net552));
 sky130_fd_sc_hd__o2111ai_1 c672 (.A1(clknet_1_1__leaf_net552),
    .A2(net549),
    .B1(net542),
    .C1(net962),
    .D1(net784),
    .Y(net553));
 sky130_fd_sc_hd__or2_1 c673 (.A(net965),
    .B(net784),
    .X(net554));
 sky130_fd_sc_hd__or4bb_1 c674 (.A(net554),
    .B(net550),
    .C_N(net547),
    .D_N(net784),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_4 c675 (.A(net705),
    .X(net556));
 sky130_fd_sc_hd__inv_4 c676 (.A(net705),
    .Y(net557));
 sky130_fd_sc_hd__or2b_1 c677 (.A(net192),
    .B_N(net72),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_1 c678 (.A(net705),
    .X(net559));
 sky130_fd_sc_hd__inv_1 c679 (.A(net761),
    .Y(net560));
 sky130_fd_sc_hd__or2_1 c68 (.A(net861),
    .B(net873),
    .X(net6));
 sky130_fd_sc_hd__inv_1 c680 (.A(net705),
    .Y(net561));
 sky130_fd_sc_hd__and2b_1 c681 (.A_N(net446),
    .B(net965),
    .X(net562));
 sky130_fd_sc_hd__or4bb_4 c682 (.A(net965),
    .B(net556),
    .C_N(net689),
    .D_N(clknet_1_1__leaf_net794),
    .X(net563));
 sky130_fd_sc_hd__or4bb_1 c683 (.A(clknet_1_0__leaf_net563),
    .B(net965),
    .C_N(net542),
    .D_N(clknet_1_1__leaf_net794),
    .X(net564));
 sky130_fd_sc_hd__or4bb_4 c684 (.A(net319),
    .B(clknet_1_1__leaf_net363),
    .C_N(net451),
    .D_N(net542),
    .X(net565));
 sky130_fd_sc_hd__nor3_1 c685 (.A(net547),
    .B(net826),
    .C(net773),
    .Y(net566));
 sky130_fd_sc_hd__mux4_4 c686 (.A0(net566),
    .A1(net562),
    .A2(clknet_1_1__leaf_net564),
    .A3(net840),
    .S0(net226),
    .S1(net952),
    .X(net567));
 sky130_fd_sc_hd__and3_2 c687 (.A(net542),
    .B(net556),
    .C(net998),
    .X(net568));
 sky130_fd_sc_hd__or4bb_2 c688 (.A(net194),
    .B(net204),
    .C_N(net568),
    .D_N(net947),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net329),
    .A1(clknet_1_0__leaf_net564),
    .A2(net327),
    .A3(net541),
    .S0(net962),
    .S1(net770),
    .X(net570));
 sky130_fd_sc_hd__and2_1 c69 (.A(net857),
    .B(net972),
    .X(net7));
 sky130_fd_sc_hd__sedfxtp_4 c690 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net363),
    .DE(net549),
    .SCD(net547),
    .SCE(net542),
    .Q(net571));
 sky130_fd_sc_hd__clkbuf_1 c691 (.A(net720),
    .X(net572));
 sky130_fd_sc_hd__or4bb_1 c692 (.A(net572),
    .B(net441),
    .C_N(net968),
    .D_N(net542),
    .X(net573));
 sky130_fd_sc_hd__mux4_4 c693 (.A0(clknet_1_0__leaf_net563),
    .A1(net226),
    .A2(net573),
    .A3(net962),
    .S0(net216),
    .S1(net766),
    .X(net574));
 sky130_fd_sc_hd__or3_2 c694 (.A(net568),
    .B(clknet_1_1__leaf_net564),
    .C(clknet_1_0__leaf_net570),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net226),
    .A1(clknet_1_0__leaf_net575),
    .A2(clknet_1_1__leaf_net570),
    .A3(net549),
    .S0(net965),
    .S1(net968),
    .X(net576));
 sky130_fd_sc_hd__or4bb_4 c696 (.A(net216),
    .B(net547),
    .C_N(net770),
    .D_N(clknet_1_0__leaf_net813),
    .X(net577));
 sky130_fd_sc_hd__or4bb_2 c697 (.A(net571),
    .B(clknet_1_0__leaf_net575),
    .C_N(net968),
    .D_N(net779),
    .X(net578));
 sky130_fd_sc_hd__a2111oi_2 c698 (.A1(net451),
    .A2(net947),
    .B1(net962),
    .C1(net770),
    .D1(clknet_1_0__leaf_net813),
    .Y(net579));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net962),
    .A1(net568),
    .A2(net826),
    .A3(net328),
    .S0(net779),
    .S1(net783),
    .X(net580));
 sky130_fd_sc_hd__nand2b_2 c70 (.A_N(net5),
    .B(net972),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net573),
    .A1(clknet_1_1__leaf_net575),
    .A2(net965),
    .A3(net580),
    .S0(net783),
    .S1(clknet_1_1__leaf_net813),
    .X(net581));
 sky130_fd_sc_hd__mux4_2 c701 (.A0(net580),
    .A1(clknet_1_0__leaf_net564),
    .A2(net573),
    .A3(net968),
    .S0(net568),
    .S1(clknet_1_0__leaf_net813),
    .X(net582));
 sky130_fd_sc_hd__mux4_2 c702 (.A0(net582),
    .A1(net562),
    .A2(net451),
    .A3(net580),
    .S0(clknet_1_0__leaf_net813),
    .S1(clknet_1_0__leaf_net814),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net580),
    .A1(clknet_1_1__leaf_net564),
    .A2(net766),
    .A3(net999),
    .S0(net779),
    .S1(net783),
    .X(net584));
 sky130_fd_sc_hd__a2111o_4 c704 (.A1(net541),
    .A2(net845),
    .B1(clknet_1_1__leaf_net584),
    .C1(net556),
    .D1(net948),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net844),
    .A1(net962),
    .A2(net204),
    .A3(clknet_1_0__leaf_net563),
    .S0(net922),
    .S1(clknet_1_1__leaf_net814),
    .X(net586));
 sky130_fd_sc_hd__mux4_4 c706 (.A0(net549),
    .A1(net543),
    .A2(net72),
    .A3(net383),
    .S0(net542),
    .S1(clknet_1_0__leaf_net812),
    .X(net587));
 sky130_fd_sc_hd__mux4_4 c707 (.A0(clknet_1_0__leaf_net563),
    .A1(net569),
    .A2(net568),
    .A3(net892),
    .S0(net328),
    .S1(net801),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net965),
    .A1(net569),
    .A2(net558),
    .A3(net556),
    .S0(net801),
    .S1(net802),
    .X(net589));
 sky130_fd_sc_hd__mux4_4 c709 (.A0(net562),
    .A1(clknet_1_1__leaf_net563),
    .A2(net840),
    .A3(net328),
    .S0(clknet_1_0__leaf_net812),
    .S1(net816),
    .X(net590));
 sky130_fd_sc_hd__o2111ai_2 c71 (.A1(net3),
    .A2(net827),
    .B1(net849),
    .C1(net873),
    .D1(net8),
    .Y(net9));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net571),
    .A1(net845),
    .A2(net892),
    .A3(net922),
    .S0(net802),
    .S1(net818),
    .X(net591));
 sky130_fd_sc_hd__mux4_2 c711 (.A0(net558),
    .A1(net962),
    .A2(clknet_1_1__leaf_net365),
    .A3(net948),
    .S0(clknet_1_1__leaf_net814),
    .S1(net815),
    .X(net592));
 sky130_fd_sc_hd__mux4_4 c712 (.A0(net592),
    .A1(net966),
    .A2(net568),
    .A3(clknet_1_1__leaf_net365),
    .S0(clknet_1_1__leaf_net814),
    .S1(net815),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net845),
    .A1(net546),
    .A2(net562),
    .A3(net569),
    .S0(net770),
    .S1(net820),
    .X(net594));
 sky130_fd_sc_hd__a2111oi_4 c714 (.A1(net542),
    .A2(net965),
    .B1(net492),
    .C1(net801),
    .D1(clknet_1_0__leaf_net814),
    .Y(net595));
 sky130_fd_sc_hd__mux4_4 c715 (.A0(clknet_1_0__leaf_net595),
    .A1(net481),
    .A2(net936),
    .A3(net801),
    .S0(net820),
    .S1(net821),
    .X(net596));
 sky130_fd_sc_hd__mux4_4 c716 (.A0(net542),
    .A1(net596),
    .A2(net541),
    .A3(net840),
    .S0(clknet_1_0__leaf_net595),
    .S1(net819),
    .X(net597));
 sky130_fd_sc_hd__o2111a_2 c717 (.A1(clknet_1_0__leaf_net595),
    .A2(net72),
    .B1(net568),
    .C1(net947),
    .D1(net820),
    .X(net598));
 sky130_fd_sc_hd__mux4_2 c718 (.A0(net947),
    .A1(net493),
    .A2(net204),
    .A3(clknet_1_0__leaf_net595),
    .S0(net815),
    .S1(net820),
    .X(net599));
 sky130_fd_sc_hd__mux4_2 c719 (.A0(clknet_1_1__leaf_net599),
    .A1(clknet_1_1__leaf_net595),
    .A2(net922),
    .A3(net816),
    .S0(net820),
    .S1(net821),
    .X(net600));
 sky130_fd_sc_hd__nor3b_1 c72 (.A(net9),
    .B(net972),
    .C_N(net879),
    .Y(net10));
 sky130_fd_sc_hd__mux4_4 c720 (.A0(net568),
    .A1(net558),
    .A2(net441),
    .A3(clknet_1_1__leaf_net595),
    .S0(net816),
    .S1(net819),
    .X(net601));
 sky130_fd_sc_hd__mux4_4 c721 (.A0(clknet_1_0__leaf_net598),
    .A1(net850),
    .A2(clknet_1_1__leaf_net595),
    .A3(net962),
    .S0(net816),
    .S1(net821),
    .X(net602));
 sky130_fd_sc_hd__mux4_4 c722 (.A0(net601),
    .A1(net597),
    .A2(clknet_1_1__leaf_net599),
    .A3(clknet_1_1__leaf_net598),
    .S0(net816),
    .S1(net821),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(clknet_1_0__leaf_net595),
    .A1(clknet_1_0__leaf_net599),
    .A2(net493),
    .A3(net481),
    .S0(net767),
    .S1(net819),
    .X(net604));
 sky130_fd_sc_hd__mux4_2 c724 (.A0(net586),
    .A1(clknet_1_1__leaf_net595),
    .A2(clknet_1_1__leaf_net599),
    .A3(clknet_1_0__leaf_net812),
    .S0(net815),
    .S1(net819),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net543),
    .A1(net483),
    .A2(clknet_1_0__leaf_net599),
    .A3(net767),
    .S0(net819),
    .S1(net821),
    .X(net606));
 sky130_fd_sc_hd__o2111ai_4 c726 (.A1(net483),
    .A2(clknet_1_1__leaf_net584),
    .B1(net952),
    .C1(net556),
    .D1(net818),
    .Y(net607));
 sky130_fd_sc_hd__o2111ai_1 c727 (.A1(net514),
    .A2(net259),
    .B1(net326),
    .C1(net803),
    .D1(net817),
    .Y(net608));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net569),
    .A1(clknet_1_1__leaf_net365),
    .A2(clknet_1_1__leaf_net399),
    .A3(clknet_1_1__leaf_net794),
    .S0(net802),
    .S1(net818),
    .X(net609));
 sky130_fd_sc_hd__sdfbbn_1 c729 (.CLK_N(clknet_4_6_0_clk),
    .D(net968),
    .RESET_B(clknet_1_1__leaf_net365),
    .SCD(clknet_1_1__leaf_net939),
    .SCE(net952),
    .SET_B(net396),
    .Q(net611),
    .Q_N(net610));
 sky130_fd_sc_hd__and2_0 c73 (.A(net837),
    .B(net873),
    .X(net11));
 sky130_fd_sc_hd__mux4_2 c730 (.A0(net571),
    .A1(clknet_1_1__leaf_net407),
    .A2(clknet_1_1__leaf_net894),
    .A3(net786),
    .S0(net804),
    .S1(net817),
    .X(net612));
 sky130_fd_sc_hd__o2111a_1 c731 (.A1(net608),
    .A2(net945),
    .B1(net610),
    .C1(net926),
    .D1(net818),
    .X(net613));
 sky130_fd_sc_hd__a2111o_4 c732 (.A1(net493),
    .A2(clknet_1_0__leaf_net399),
    .B1(net804),
    .C1(clknet_1_1__leaf_net812),
    .D1(net817),
    .X(net940));
 sky130_fd_sc_hd__mux4_4 c733 (.A0(net556),
    .A1(clknet_1_0__leaf_net940),
    .A2(net934),
    .A3(net906),
    .S0(clknet_1_1__leaf_net812),
    .S1(net817),
    .X(net614));
 sky130_fd_sc_hd__o2111a_2 c734 (.A1(clknet_1_1__leaf_net517),
    .A2(net840),
    .B1(clknet_1_0__leaf_net940),
    .C1(net892),
    .D1(net818),
    .X(net615));
 sky130_fd_sc_hd__mux4_4 c735 (.A0(clknet_1_1__leaf_net407),
    .A1(net613),
    .A2(net840),
    .A3(clknet_1_1__leaf_net517),
    .S0(clknet_1_0__leaf_net940),
    .S1(net906),
    .X(net616));
 sky130_fd_sc_hd__a2111oi_1 c736 (.A1(net571),
    .A2(clknet_1_0__leaf_net940),
    .B1(net783),
    .C1(net786),
    .D1(net818),
    .Y(net617));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net556),
    .A1(net617),
    .A2(net571),
    .A3(clknet_1_0__leaf_net940),
    .S0(net518),
    .S1(clknet_1_1__leaf_net812),
    .X(net618));
 sky130_fd_sc_hd__sdfbbp_1 c738 (.CLK(clknet_4_7_0_clk),
    .D(net614),
    .RESET_B(net612),
    .SCD(clknet_1_1__leaf_net517),
    .SCE(net968),
    .SET_B(net785),
    .Q(net890),
    .Q_N(net619));
 sky130_fd_sc_hd__o2111ai_4 c739 (.A1(net546),
    .A2(net890),
    .B1(net945),
    .C1(net906),
    .D1(net817),
    .Y(net620));
 sky130_fd_sc_hd__or2b_1 c74 (.A(net4),
    .B_N(net8),
    .X(net12));
 sky130_fd_sc_hd__o2111ai_1 c740 (.A1(net493),
    .A2(net620),
    .B1(net890),
    .C1(net571),
    .D1(clknet_1_1__leaf_net794),
    .Y(net621));
 sky130_fd_sc_hd__mux4_2 c741 (.A0(net259),
    .A1(clknet_1_1__leaf_net940),
    .A2(net934),
    .A3(net782),
    .S0(net784),
    .S1(net906),
    .X(net622));
 sky130_fd_sc_hd__mux4_2 c742 (.A0(net618),
    .A1(net569),
    .A2(net619),
    .A3(net875),
    .S0(net620),
    .S1(net755),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net556),
    .A1(net620),
    .A2(net952),
    .A3(clknet_1_1__leaf_net940),
    .S0(net784),
    .S1(net785),
    .X(net624));
 sky130_fd_sc_hd__mux4_4 c744 (.A0(net620),
    .A1(net556),
    .A2(net235),
    .A3(net769),
    .S0(net803),
    .S1(net971),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net259),
    .A1(net329),
    .A2(net620),
    .A3(clknet_1_1__leaf_net407),
    .S0(net926),
    .S1(net823),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net556),
    .A1(net483),
    .A2(net619),
    .A3(net926),
    .S0(net770),
    .S1(net823),
    .X(net627));
 sky130_fd_sc_hd__o2111a_1 c747 (.A1(net235),
    .A2(net769),
    .B1(net784),
    .C1(net817),
    .D1(net823),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net1009),
    .A1(net898),
    .A2(clknet_1_1__leaf_net939),
    .A3(net796),
    .S0(net808),
    .S1(net971),
    .X(net629));
 sky130_fd_sc_hd__mux4_4 c749 (.A0(net627),
    .A1(net888),
    .A2(net886),
    .A3(net810),
    .S0(net811),
    .S1(net822),
    .X(net630));
 sky130_fd_sc_hd__and2b_1 c75 (.A_N(net7),
    .B(net972),
    .X(net13));
 sky130_fd_sc_hd__mux4_2 c750 (.A0(net327),
    .A1(clknet_1_0__leaf_net395),
    .A2(net886),
    .A3(clknet_1_1__leaf_net940),
    .S0(net792),
    .S1(net971),
    .X(net631));
 sky130_fd_sc_hd__mux4_4 c751 (.A0(net497),
    .A1(net538),
    .A2(net327),
    .A3(net838),
    .S0(clknet_1_0__leaf_net584),
    .S1(net875),
    .X(net632));
 sky130_fd_sc_hd__mux4_2 c752 (.A0(net630),
    .A1(net622),
    .A2(clknet_1_1__leaf_net939),
    .A3(net892),
    .S0(net802),
    .S1(net822),
    .X(net633));
 sky130_fd_sc_hd__mux4_2 c753 (.A0(net329),
    .A1(net1009),
    .A2(net496),
    .A3(net783),
    .S0(net802),
    .S1(net807),
    .X(net634));
 sky130_fd_sc_hd__mux4_2 c754 (.A0(net611),
    .A1(net634),
    .A2(clknet_1_0__leaf_net584),
    .A3(clknet_1_1__leaf_net894),
    .S0(net783),
    .S1(net792),
    .X(net635));
 sky130_fd_sc_hd__mux4_2 c755 (.A0(net631),
    .A1(clknet_1_0__leaf_net584),
    .A2(net952),
    .A3(net350),
    .S0(net634),
    .S1(net778),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net82),
    .A1(net634),
    .A2(net774),
    .A3(net778),
    .S0(net782),
    .S1(net971),
    .X(net637));
 sky130_fd_sc_hd__mux4_4 c757 (.A0(net987),
    .A1(clknet_1_1__leaf_net940),
    .A2(net875),
    .A3(net888),
    .S0(net971),
    .S1(net823),
    .X(net638));
 sky130_fd_sc_hd__mux4_4 c758 (.A0(net634),
    .A1(net755),
    .A2(net796),
    .A3(net811),
    .S0(net971),
    .S1(net823),
    .X(net639));
 sky130_fd_sc_hd__mux4_2 c759 (.A0(net637),
    .A1(net540),
    .A2(net952),
    .A3(net634),
    .S0(net810),
    .S1(net811),
    .X(net640));
 sky130_fd_sc_hd__or2_1 c76 (.A(net13),
    .B(net972),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net950),
    .A1(net634),
    .A2(net497),
    .A3(net611),
    .S0(net802),
    .S1(net971),
    .X(net641));
 sky130_fd_sc_hd__mux4_4 c761 (.A0(clknet_1_1__leaf_net395),
    .A1(clknet_1_1__leaf_net638),
    .A2(net634),
    .A3(net82),
    .S0(net768),
    .S1(net792),
    .X(net642));
 sky130_fd_sc_hd__mux4_2 c762 (.A0(net519),
    .A1(clknet_1_0__leaf_net638),
    .A2(net497),
    .A3(net875),
    .S0(net935),
    .S1(net971),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net628),
    .A1(clknet_1_1__leaf_net584),
    .A2(net875),
    .A3(net634),
    .S0(net778),
    .S1(net810),
    .X(net644));
 sky130_fd_sc_hd__mux4_2 c764 (.A0(net888),
    .A1(clknet_1_1__leaf_net643),
    .A2(net634),
    .A3(clknet_1_1__leaf_net939),
    .S0(net810),
    .S1(net822),
    .X(net645));
 sky130_fd_sc_hd__mux4_2 c765 (.A0(net350),
    .A1(net524),
    .A2(net887),
    .A3(net792),
    .S0(net935),
    .S1(net895),
    .X(net646));
 sky130_fd_sc_hd__mux4_2 c766 (.A0(net386),
    .A1(net639),
    .A2(net634),
    .A3(clknet_1_0__leaf_net584),
    .S0(net971),
    .S1(net895),
    .X(net647));
 sky130_fd_sc_hd__mux4_2 c767 (.A0(clknet_1_0__leaf_net643),
    .A1(net887),
    .A2(net781),
    .A3(net782),
    .S0(net792),
    .S1(net895),
    .X(net648));
 sky130_fd_sc_hd__mux4_4 c768 (.A0(net641),
    .A1(net640),
    .A2(net936),
    .A3(net781),
    .S0(net971),
    .S1(net895),
    .X(net649));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net642),
    .A1(net649),
    .A2(net768),
    .A3(net781),
    .S0(net811),
    .S1(net895),
    .X(net650));
 sky130_fd_sc_hd__or2_1 c77 (.A(net6),
    .B(net14),
    .X(net15));
 sky130_fd_sc_hd__and2b_1 c78 (.A_N(net10),
    .B(net972),
    .X(net16));
 sky130_fd_sc_hd__and2b_1 c79 (.A_N(net16),
    .B(net11),
    .X(net17));
 sky130_fd_sc_hd__nand3b_4 c80 (.A_N(net849),
    .B(net972),
    .C(net961),
    .Y(net18));
 sky130_fd_sc_hd__mux4_2 c81 (.A0(net11),
    .A1(net1),
    .A2(net17),
    .A3(net7),
    .S0(net846),
    .S1(net842),
    .X(net19));
 sky130_fd_sc_hd__nor3b_1 c82 (.A(net17),
    .B(net9),
    .C_N(net961),
    .Y(net20));
 sky130_fd_sc_hd__nand3_1 c83 (.A(net18),
    .B(net959),
    .C(net961),
    .Y(net21));
 sky130_fd_sc_hd__or2b_1 c84 (.A(net12),
    .B_N(net861),
    .X(net22));
 sky130_fd_sc_hd__or2_4 c85 (.A(net863),
    .B(net3),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 c86 (.A0(net22),
    .A1(net7),
    .A2(net23),
    .A3(net842),
    .S0(net13),
    .S1(net846),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 c87 (.A0(net24),
    .A1(net5),
    .A2(net14),
    .A3(net18),
    .S0(net875),
    .S1(net873),
    .X(net25));
 sky130_fd_sc_hd__nand2b_1 c88 (.A_N(net25),
    .B(net24),
    .Y(net26));
 sky130_fd_sc_hd__or2_1 c89 (.A(net846),
    .B(net871),
    .X(net27));
 sky130_fd_sc_hd__nor2_2 c90 (.A(net26),
    .B(net870),
    .Y(net28));
 sky130_fd_sc_hd__and2_2 c91 (.A(net835),
    .B(net18),
    .X(net29));
 sky130_fd_sc_hd__nor3b_4 c92 (.A(net859),
    .B(net28),
    .C_N(net972),
    .Y(net30));
 sky130_fd_sc_hd__or4bb_4 c93 (.A(net865),
    .B(net29),
    .C_N(net957),
    .D_N(net961),
    .X(net923));
 sky130_fd_sc_hd__or2_4 c94 (.A(net866),
    .B(net29),
    .X(net31));
 sky130_fd_sc_hd__and2_1 c95 (.A(net24),
    .B(net26),
    .X(net909));
 sky130_fd_sc_hd__and2_1 c96 (.A(net27),
    .B(net877),
    .X(net32));
 sky130_fd_sc_hd__nand2_1 c97 (.A(net868),
    .B(net31),
    .Y(net33));
 sky130_fd_sc_hd__and3b_1 c98 (.A_N(net30),
    .B(net28),
    .C(net958),
    .X(net34));
 sky130_fd_sc_hd__nor2_2 c99 (.A(net33),
    .B(net958),
    .Y(net35));
 sky130_fd_sc_hd__a2111o_1 merge790 (.A1(net341),
    .A2(net320),
    .B1(net322),
    .C1(net77),
    .D1(net1011),
    .X(net651));
 sky130_fd_sc_hd__mux4_2 merge791 (.A0(clknet_1_0__leaf_net425),
    .A1(clknet_1_1__leaf_net292),
    .A2(net350),
    .A3(clknet_1_0__leaf_net423),
    .S0(clknet_1_1__leaf_net289),
    .S1(net31),
    .X(net652));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net112),
    .A1(net116),
    .A2(net204),
    .A3(net236),
    .S0(net945),
    .S1(net722),
    .X(net653));
 sky130_fd_sc_hd__or4bb_1 merge793 (.A(net434),
    .B(net319),
    .C_N(net197),
    .D_N(net322),
    .X(net654));
 sky130_fd_sc_hd__mux4_2 merge794 (.A0(net157),
    .A1(clknet_1_1__leaf_net169),
    .A2(net55),
    .A3(net176),
    .S0(net173),
    .S1(net694),
    .X(net655));
 sky130_fd_sc_hd__o2111a_4 merge795 (.A1(clknet_1_0__leaf_net439),
    .A2(net435),
    .B1(net200),
    .C1(net941),
    .D1(net948),
    .X(net656));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net449),
    .A1(net451),
    .A2(net344),
    .A3(net857),
    .S0(net950),
    .S1(net319),
    .X(net657));
 sky130_fd_sc_hd__a2111o_4 merge797 (.A1(clknet_1_1__leaf_net135),
    .A2(net157),
    .B1(clknet_1_1__leaf_net140),
    .C1(net19),
    .D1(clknet_1_0__leaf_net161),
    .X(net658));
 sky130_fd_sc_hd__o2111ai_1 merge798 (.A1(net119),
    .A2(net875),
    .B1(net879),
    .C1(net857),
    .D1(net128),
    .Y(net659));
 sky130_fd_sc_hd__or4bb_4 merge799 (.A(net953),
    .B(net236),
    .C_N(clknet_1_0__leaf_net372),
    .D_N(net126),
    .X(net660));
 sky130_fd_sc_hd__or4bb_1 merge800 (.A(net223),
    .B(net233),
    .C_N(net335),
    .D_N(net340),
    .X(net661));
 sky130_fd_sc_hd__o2111a_2 merge801 (.A1(net242),
    .A2(clknet_1_0__leaf_net160),
    .B1(net960),
    .C1(net279),
    .D1(net270),
    .X(net662));
 sky130_fd_sc_hd__mux4_1 merge802 (.A0(net214),
    .A1(net833),
    .A2(net942),
    .A3(net842),
    .S0(net851),
    .S1(net216),
    .X(net663));
 sky130_fd_sc_hd__or4bb_1 merge803 (.A(net351),
    .B(net319),
    .C_N(net233),
    .D_N(net349),
    .X(net664));
 sky130_fd_sc_hd__mux4_2 merge804 (.A0(net91),
    .A1(clknet_1_0__leaf_net145),
    .A2(clknet_1_0__leaf_net146),
    .A3(net114),
    .S0(clknet_1_0__leaf_net135),
    .S1(net19),
    .X(net665));
 sky130_fd_sc_hd__mux4_2 merge805 (.A0(net872),
    .A1(net119),
    .A2(net8),
    .A3(net223),
    .S0(net95),
    .S1(net216),
    .X(net666));
 sky130_fd_sc_hd__mux4_4 merge806 (.A0(net121),
    .A1(net879),
    .A2(net961),
    .A3(clknet_1_0__leaf_net148),
    .S0(net183),
    .S1(net919),
    .X(net667));
 sky130_fd_sc_hd__mux4_4 merge807 (.A0(net236),
    .A1(net269),
    .A2(net386),
    .A3(clknet_1_0__leaf_net292),
    .S0(net966),
    .S1(net261),
    .X(net668));
 sky130_fd_sc_hd__mux4_1 merge808 (.A0(net421),
    .A1(clknet_1_0__leaf_net254),
    .A2(net30),
    .A3(net411),
    .S0(net122),
    .S1(net741),
    .X(net669));
 sky130_fd_sc_hd__mux4_2 merge809 (.A0(net218),
    .A1(net116),
    .A2(net238),
    .A3(net23),
    .S0(clknet_1_0__leaf_net160),
    .S1(net162),
    .X(net670));
 sky130_fd_sc_hd__mux4_4 merge810 (.A0(net411),
    .A1(net410),
    .A2(net386),
    .A3(clknet_1_1__leaf_net254),
    .S0(net897),
    .S1(net383),
    .X(net671));
 sky130_fd_sc_hd__mux4_1 merge811 (.A0(net463),
    .A1(net459),
    .A2(net464),
    .A3(clknet_1_0__leaf_net570),
    .S0(net216),
    .S1(net226),
    .X(net672));
 sky130_fd_sc_hd__mux4_4 merge812 (.A0(net942),
    .A1(net216),
    .A2(net995),
    .A3(net376),
    .S0(net370),
    .S1(net907),
    .X(net673));
 sky130_fd_sc_hd__a2111o_1 merge813 (.A1(clknet_1_1__leaf_net438),
    .A2(net847),
    .B1(net555),
    .C1(net446),
    .D1(clknet_1_0__leaf_net552),
    .X(net674));
 sky130_fd_sc_hd__mux4_2 merge814 (.A0(clknet_1_0__leaf_net438),
    .A1(net900),
    .A2(net432),
    .A3(net247),
    .S0(net243),
    .S1(net244),
    .X(net675));
 sky130_fd_sc_hd__mux4_1 merge815 (.A0(net231),
    .A1(net942),
    .A2(net216),
    .A3(net342),
    .S0(net349),
    .S1(net1020),
    .X(net676));
 sky130_fd_sc_hd__mux4_4 merge816 (.A0(net114),
    .A1(net91),
    .A2(net873),
    .A3(net239),
    .S0(net241),
    .S1(net243),
    .X(net677));
 sky130_fd_sc_hd__mux4_1 merge817 (.A0(net428),
    .A1(net431),
    .A2(net941),
    .A3(net432),
    .S0(net434),
    .S1(net326),
    .X(net678));
 sky130_fd_sc_hd__mux4_4 merge818 (.A0(net433),
    .A1(net431),
    .A2(net427),
    .A3(clknet_1_0__leaf_net442),
    .S0(clknet_1_0__leaf_net447),
    .S1(net943),
    .X(net679));
 sky130_fd_sc_hd__mux4_1 merge819 (.A0(net431),
    .A1(net435),
    .A2(net339),
    .A3(net322),
    .S0(clknet_1_0__leaf_net438),
    .S1(net965),
    .X(net680));
 sky130_fd_sc_hd__dfrbp_1 merge820 (.CLK(clknet_4_2_0_clk),
    .D(net380),
    .RESET_B(net660),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dfrbp_1 merge821 (.CLK(clknet_4_1_0_clk),
    .D(net458),
    .RESET_B(net470),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__dfrtn_1 merge822 (.CLK_N(clknet_4_4_0_clk),
    .D(net444),
    .RESET_B(net656),
    .Q(net685));
 sky130_fd_sc_hd__dfrtp_2 merge823 (.CLK(clknet_4_0_0_clk),
    .D(net333),
    .RESET_B(net651),
    .Q(net686));
 sky130_fd_sc_hd__or2_1 merge824 (.A(net607),
    .B(net609),
    .X(net687));
 sky130_fd_sc_hd__dfrtp_4 merge825 (.CLK(clknet_4_3_0_clk),
    .D(net474),
    .RESET_B(net485),
    .Q(net903));
 sky130_fd_sc_hd__and2b_4 merge826 (.A_N(net567),
    .B(net578),
    .X(net688));
 sky130_fd_sc_hd__dfrtp_1 merge827 (.CLK(clknet_4_0_0_clk),
    .RESET_B(net103),
    .Q(net104));
 sky130_fd_sc_hd__nand2_1 merge828 (.A(net266),
    .B(net277),
    .Y(net690));
 sky130_fd_sc_hd__nand2_2 merge829 (.A(net298),
    .B(net304),
    .Y(net691));
 sky130_fd_sc_hd__nand2_1 merge830 (.A(net677),
    .B(net127),
    .Y(net692));
 sky130_fd_sc_hd__dfsbp_2 merge831 (.CLK(clknet_4_10_0_clk),
    .D(net62),
    .SET_B(net61),
    .Q(net694),
    .Q_N(net693));
 sky130_fd_sc_hd__nand2_1 merge832 (.A(net245),
    .B(net246),
    .Y(net695));
 sky130_fd_sc_hd__or2_2 merge833 (.A(net505),
    .B(net498),
    .X(net696));
 sky130_fd_sc_hd__nand2b_2 merge834 (.A_N(net168),
    .B(net167),
    .Y(net697));
 sky130_fd_sc_hd__or2_1 merge835 (.A(net181),
    .B(net184),
    .X(net698));
 sky130_fd_sc_hd__dfsbp_1 merge836 (.CLK(clknet_4_12_0_clk),
    .D(net397),
    .SET_B(net398),
    .Q(net700),
    .Q_N(net699));
 sky130_fd_sc_hd__nor2b_2 merge837 (.A(net650),
    .B_N(net629),
    .Y(net701));
 sky130_fd_sc_hd__nor2_2 merge838 (.A(net408),
    .B(net418),
    .Y(net702));
 sky130_fd_sc_hd__nand2_2 merge839 (.A(net585),
    .B(net587),
    .Y(net703));
 sky130_fd_sc_hd__dfstp_2 merge840 (.CLK(clknet_4_8_0_clk),
    .D(net659),
    .SET_B(net665),
    .Q(net704));
 sky130_fd_sc_hd__dfstp_1 merge841 (.CLK(clknet_4_4_0_clk),
    .D(net654),
    .SET_B(net674),
    .Q(net705));
 sky130_fd_sc_hd__nand2b_1 merge842 (.A_N(net362),
    .B(net360),
    .Y(net706));
 sky130_fd_sc_hd__or2_4 merge843 (.A(net528),
    .B(net529),
    .X(net707));
 sky130_fd_sc_hd__nor2_2 merge844 (.A(net281),
    .B(net285),
    .Y(net708));
 sky130_fd_sc_hd__and2b_1 merge845 (.A_N(net663),
    .B(net673),
    .X(net709));
 sky130_fd_sc_hd__nor2b_1 merge846 (.A(net701),
    .B_N(net615),
    .Y(net710));
 sky130_fd_sc_hd__nor2_1 merge847 (.A(net583),
    .B(net661),
    .Y(net711));
 sky130_fd_sc_hd__and2b_2 merge848 (.A_N(net253),
    .B(net295),
    .X(net712));
 sky130_fd_sc_hd__or2b_4 merge849 (.A(net426),
    .B_N(net318),
    .X(net713));
 sky130_fd_sc_hd__nor2b_2 merge850 (.A(net189),
    .B_N(net317),
    .Y(net714));
 sky130_fd_sc_hd__and2b_1 merge851 (.A_N(net187),
    .B(net666),
    .X(net715));
 sky130_fd_sc_hd__nand2_1 merge852 (.A(net305),
    .B(net315),
    .Y(net716));
 sky130_fd_sc_hd__dfstp_4 merge853 (.CLK(clknet_4_0_0_clk),
    .D(net664),
    .SET_B(net676),
    .Q(net717));
 sky130_fd_sc_hd__nor2b_4 merge854 (.A(net537),
    .B_N(net312),
    .Y(net718));
 sky130_fd_sc_hd__nand2b_4 merge855 (.A_N(net591),
    .B(net648),
    .Y(net719));
 sky130_fd_sc_hd__dlrbn_1 merge856 (.D(net706),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net672),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dlrbn_1 merge857 (.D(net709),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net220),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__nor2_1 merge858 (.A(net539),
    .B(net718),
    .Y(net724));
 sky130_fd_sc_hd__or2b_1 merge859 (.A(net633),
    .B_N(net646),
    .X(net725));
 sky130_fd_sc_hd__or2b_4 merge860 (.A(net250),
    .B_N(net255),
    .X(net726));
 sky130_fd_sc_hd__dlrbp_1 merge861 (.D(net708),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net671),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__nor2b_1 merge862 (.A(net311),
    .B_N(net713),
    .Y(net729));
 sky130_fd_sc_hd__nor2b_4 merge863 (.A(net670),
    .B_N(net521),
    .Y(net730));
 sky130_fd_sc_hd__or2b_1 merge864 (.A(net626),
    .B_N(net624),
    .X(net731));
 sky130_fd_sc_hd__dlrbp_1 merge865 (.D(net712),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net695),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__dlrtn_4 merge866 (.D(net667),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net144),
    .Q(net734));
 sky130_fd_sc_hd__dlrtn_2 merge867 (.D(net653),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net668),
    .Q(net735));
 sky130_fd_sc_hd__and2_1 merge868 (.A(net635),
    .B(net636),
    .X(net736));
 sky130_fd_sc_hd__nand2_2 merge869 (.A(net272),
    .B(net275),
    .Y(net737));
 sky130_fd_sc_hd__nor2b_1 merge870 (.A(net588),
    .B_N(net623),
    .Y(net738));
 sky130_fd_sc_hd__dlrtn_1 merge871 (.D(net731),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net687),
    .Q(net926));
 sky130_fd_sc_hd__nor2_2 merge872 (.A(net600),
    .B(net606),
    .Y(net739));
 sky130_fd_sc_hd__dlrtp_1 merge873 (.D(net655),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net716),
    .Q(net740));
 sky130_fd_sc_hd__dlrtp_4 merge874 (.D(net658),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net697),
    .Q(net741));
 sky130_fd_sc_hd__dlrtp_2 merge875 (.D(net185),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net698),
    .Q(net919));
 sky130_fd_sc_hd__edfxbp_1 merge876 (.CLK(clknet_4_2_0_clk),
    .D(net692),
    .DE(net118),
    .Q(net743),
    .Q_N(net742));
 sky130_fd_sc_hd__or2_2 merge877 (.A(net602),
    .B(net605),
    .X(net744));
 sky130_fd_sc_hd__edfxtp_1 merge878 (.CLK(clknet_4_6_0_clk),
    .D(net491),
    .DE(net487),
    .Q(net913));
 sky130_fd_sc_hd__and2_2 merge879 (.A(net604),
    .B(net736),
    .X(net745));
 sky130_fd_sc_hd__sdlclkp_1 merge880 (.CLK(clknet_4_1_0_clk),
    .GATE(net675),
    .SCE(net678),
    .GCLK(net746));
 sky130_fd_sc_hd__sdlclkp_2 merge881 (.CLK(clknet_4_9_0_clk),
    .GATE(net690),
    .SCE(net274),
    .GCLK(net747));
 sky130_fd_sc_hd__sdlclkp_4 merge882 (.CLK(clknet_4_11_0_clk),
    .GATE(net702),
    .SCE(net669),
    .GCLK(net748));
 sky130_fd_sc_hd__dfrbp_1 merge883 (.CLK(clknet_4_11_0_clk),
    .D(net662),
    .RESET_B(net691),
    .Q(net750),
    .Q_N(net749));
 sky130_fd_sc_hd__dfrbp_1 merge884 (.CLK(clknet_4_0_0_clk),
    .D(net323),
    .RESET_B(net385),
    .Q(net752),
    .Q_N(net751));
 sky130_fd_sc_hd__dfrtn_1 merge885 (.CLK_N(clknet_4_14_0_clk),
    .D(net420),
    .RESET_B(net316),
    .Q(net753));
 sky130_fd_sc_hd__dfrtp_4 merge886 (.CLK(clknet_4_9_0_clk),
    .D(net703),
    .RESET_B(net314),
    .Q(net934));
 sky130_fd_sc_hd__dfrtp_4 merge887 (.CLK(clknet_4_14_0_clk),
    .D(net719),
    .RESET_B(net301),
    .Q(net936));
 sky130_fd_sc_hd__dfrtp_4 merge888 (.CLK(clknet_4_11_0_clk),
    .D(net499),
    .RESET_B(net313),
    .Q(net754));
 sky130_fd_sc_hd__dfsbp_1 merge889 (.CLK(clknet_4_6_0_clk),
    .D(net486),
    .SET_B(net710),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__or2_2 merge890 (.A(net282),
    .B(net303),
    .X(net757));
 sky130_fd_sc_hd__dfsbp_1 merge891 (.CLK(clknet_4_11_0_clk),
    .D(net417),
    .SET_B(net714),
    .Q(net759),
    .Q_N(net758));
 sky130_fd_sc_hd__dfstp_2 merge892 (.CLK(clknet_4_12_0_clk),
    .D(net401),
    .SET_B(net369),
    .Q(net911));
 sky130_fd_sc_hd__dfstp_2 merge893 (.CLK(clknet_4_12_0_clk),
    .D(net507),
    .SET_B(net707),
    .Q(net760));
 sky130_fd_sc_hd__dfstp_1 merge894 (.CLK(clknet_4_4_0_clk),
    .D(net679),
    .SET_B(net680),
    .Q(net761));
 sky130_fd_sc_hd__dlrbn_2 merge895 (.D(net726),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net730),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__dlrbn_1 merge896 (.D(net657),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net520),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__dlrbp_1 merge897 (.D(net744),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net688),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__dlrbp_1 merge898 (.D(net739),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net725),
    .Q(net769),
    .Q_N(net768));
 sky130_fd_sc_hd__dlrtn_2 merge899 (.D(net738),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net565),
    .Q(net770));
 sky130_fd_sc_hd__dlrtn_1 merge900 (.D(net287),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net294));
 sky130_fd_sc_hd__dlrtn_2 merge901 (.D(net374),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net336),
    .Q(net771));
 sky130_fd_sc_hd__dlrtp_1 merge902 (.D(net533),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net652),
    .Q(net772));
 sky130_fd_sc_hd__dlrtp_4 merge903 (.D(net456),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net711),
    .Q(net773));
 sky130_fd_sc_hd__dlrtp_4 merge904 (.D(net461),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net724),
    .Q(net774));
 sky130_fd_sc_hd__edfxbp_1 merge905 (.CLK(clknet_4_14_0_clk),
    .D(net484),
    .DE(net307),
    .Q(net775),
    .Q_N(net889));
 sky130_fd_sc_hd__edfxtp_1 merge906 (.CLK(clknet_4_13_0_clk),
    .D(net469),
    .DE(net644),
    .Q(net887));
 sky130_fd_sc_hd__sdlclkp_1 merge907 (.CLK(clknet_4_10_0_clk),
    .GATE(net715),
    .SCE(net190),
    .GCLK(net776));
 sky130_fd_sc_hd__sdlclkp_2 merge908 (.CLK(clknet_4_8_0_clk),
    .GATE(net737),
    .SCE(net757),
    .GCLK(net777));
 sky130_fd_sc_hd__sdlclkp_4 merge909 (.CLK(clknet_4_10_0_clk),
    .GATE(net729),
    .SCE(net177),
    .GCLK(net901));
 sky130_fd_sc_hd__dfrbp_2 merge910 (.CLK(clknet_4_7_0_clk),
    .D(net577),
    .RESET_B(net632),
    .Q(net779),
    .Q_N(net778));
 sky130_fd_sc_hd__dfrbp_1 merge911 (.CLK(clknet_4_13_0_clk),
    .D(net647),
    .RESET_B(net400),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dfrtn_1 merge912 (.CLK_N(clknet_4_4_0_clk),
    .D(net462),
    .RESET_B(net745),
    .Q(net782));
 sky130_fd_sc_hd__dfrtp_4 merge913 (.CLK(clknet_4_6_0_clk),
    .D(net579),
    .RESET_B(net508),
    .Q(net783));
 sky130_fd_sc_hd__dfrtp_4 merge914 (.CLK(clknet_4_4_0_clk),
    .D(net553),
    .RESET_B(net384),
    .Q(net922));
 sky130_fd_sc_hd__dfrtp_4 merge915 (.CLK(clknet_4_5_0_clk),
    .D(net551),
    .RESET_B(net621),
    .Q(net784));
 sky130_fd_sc_hd__dfsbp_1 merge916 (.CLK(clknet_4_13_0_clk),
    .D(net696),
    .SET_B(net616),
    .Q(net786),
    .Q_N(net785));
 sky130_fd_sc_hd__dfxbp_1 s917 (.CLK(clknet_4_2_0_clk),
    .D(net125),
    .Q(net788),
    .Q_N(net787));
 sky130_fd_sc_hd__dfxbp_1 s918 (.CLK(clknet_4_10_0_clk),
    .D(net171),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dfxtp_2 s919 (.CLK(clknet_4_9_0_clk),
    .D(net273),
    .Q(net791));
 sky130_fd_sc_hd__dfxtp_4 s920 (.CLK(clknet_4_14_0_clk),
    .D(net296),
    .Q(net792));
 sky130_fd_sc_hd__dfxtp_4 s921 (.CLK(clknet_4_11_0_clk),
    .D(net310),
    .Q(net793));
 sky130_fd_sc_hd__dlclkp_1 s922 (.CLK(clknet_4_1_0_clk),
    .GATE(net352),
    .GCLK(net794));
 sky130_fd_sc_hd__dlclkp_2 s923 (.CLK(clknet_4_12_0_clk),
    .GATE(net405),
    .GCLK(net795));
 sky130_fd_sc_hd__dlclkp_4 s924 (.CLK(clknet_4_14_0_clk),
    .GATE(net415),
    .GCLK(net904));
 sky130_fd_sc_hd__dlxbn_2 s925 (.D(net424),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net935),
    .Q_N(net796));
 sky130_fd_sc_hd__dlxbn_1 s926 (.D(net468),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net798),
    .Q_N(net797));
 sky130_fd_sc_hd__dlxbp_1 s927 (.D(net471),
    .GATE(clknet_4_4_0_clk),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dlxtn_4 s928 (.D(net490),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net906));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net494),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net801));
 sky130_fd_sc_hd__dlxtn_4 s930 (.D(net495),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net802));
 sky130_fd_sc_hd__dlxtp_1 s931 (.D(net501),
    .GATE(clknet_4_12_0_clk),
    .Q(net803));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s932 (.D(net506),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net804));
 sky130_fd_sc_hd__dfxbp_1 s933 (.CLK(clknet_4_15_0_clk),
    .D(net525),
    .Q(net806),
    .Q_N(net805));
 sky130_fd_sc_hd__dfxbp_2 s934 (.CLK(clknet_4_15_0_clk),
    .D(net526),
    .Q(net808),
    .Q_N(net807));
 sky130_fd_sc_hd__dfxtp_1 s935 (.CLK(clknet_4_15_0_clk),
    .D(net530),
    .Q(net809));
 sky130_fd_sc_hd__dfxtp_4 s936 (.CLK(clknet_4_15_0_clk),
    .D(net531),
    .Q(net810));
 sky130_fd_sc_hd__dfxtp_1 s937 (.CLK(clknet_4_15_0_clk),
    .D(net532),
    .Q(net811));
 sky130_fd_sc_hd__dlclkp_1 s938 (.CLK(clknet_4_5_0_clk),
    .GATE(net574),
    .GCLK(net812));
 sky130_fd_sc_hd__dlclkp_2 s939 (.CLK(clknet_4_5_0_clk),
    .GATE(net576),
    .GCLK(net813));
 sky130_fd_sc_hd__dlclkp_4 s940 (.CLK(clknet_4_5_0_clk),
    .GATE(net581),
    .GCLK(net814));
 sky130_fd_sc_hd__dlxbn_2 s941 (.D(net589),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net816),
    .Q_N(net815));
 sky130_fd_sc_hd__dlxbn_2 s942 (.D(net590),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net818),
    .Q_N(net817));
 sky130_fd_sc_hd__dlxbp_1 s943 (.D(net593),
    .GATE(clknet_4_5_0_clk),
    .Q(net820),
    .Q_N(net819));
 sky130_fd_sc_hd__dlxtn_1 s944 (.D(net594),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net821));
 sky130_fd_sc_hd__dlxtn_1 s945 (.D(net603),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net822));
 sky130_fd_sc_hd__dlxtn_1 s946 (.D(net625),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net823));
 sky130_fd_sc_hd__dlxtp_1 s947 (.D(net645),
    .GATE(clknet_4_15_0_clk),
    .Q(net895));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net824));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_8 input3 (.A(in10),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net827));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(in12),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(in13),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net830));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net831));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(in17),
    .X(net833));
 sky130_fd_sc_hd__buf_1 input11 (.A(in18),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(in19),
    .X(net835));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net836));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net838));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net839));
 sky130_fd_sc_hd__buf_4 input17 (.A(in23),
    .X(net840));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net841));
 sky130_fd_sc_hd__buf_2 input19 (.A(in25),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in26),
    .X(net843));
 sky130_fd_sc_hd__buf_4 input21 (.A(in27),
    .X(net844));
 sky130_fd_sc_hd__buf_2 input22 (.A(in28),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(in29),
    .X(net846));
 sky130_fd_sc_hd__buf_2 input24 (.A(in3),
    .X(net847));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(in30),
    .X(net848));
 sky130_fd_sc_hd__buf_1 input26 (.A(in31),
    .X(net849));
 sky130_fd_sc_hd__buf_4 input27 (.A(in32),
    .X(net850));
 sky130_fd_sc_hd__buf_2 input28 (.A(in33),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(in34),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(in35),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net854));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net855));
 sky130_fd_sc_hd__buf_1 input33 (.A(in38),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(in39),
    .X(net857));
 sky130_fd_sc_hd__buf_1 input35 (.A(in4),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(in40),
    .X(net859));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net860));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net861));
 sky130_fd_sc_hd__buf_4 input39 (.A(in43),
    .X(net862));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net863));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(in46),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(in47),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in49),
    .X(net868));
 sky130_fd_sc_hd__buf_4 input46 (.A(in5),
    .X(net869));
 sky130_fd_sc_hd__buf_2 input47 (.A(in50),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(in51),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(in52),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net873));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(in54),
    .X(net874));
 sky130_fd_sc_hd__buf_4 input52 (.A(in55),
    .X(net875));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in57),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(in58),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net879));
 sky130_fd_sc_hd__buf_1 input57 (.A(in6),
    .X(net880));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(in60),
    .X(net881));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net882));
 sky130_fd_sc_hd__buf_1 input60 (.A(in7),
    .X(net883));
 sky130_fd_sc_hd__buf_1 input61 (.A(in8),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(in9),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net886),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net887),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net888),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net889),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net890),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output68 (.A(net891),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net892),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net893),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(clknet_1_0__leaf_net894),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net895),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output73 (.A(net948),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output74 (.A(net897),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output75 (.A(net898),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(clknet_1_1__leaf_net899),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output77 (.A(net900),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(clknet_1_1__leaf_net901),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output79 (.A(net902),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net903),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(clknet_1_1__leaf_net904),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(clknet_1_1__leaf_net905),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net906),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output84 (.A(net907),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output85 (.A(net908),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output86 (.A(net958),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_1__leaf_net910),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output88 (.A(net911),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net978),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net913),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net914),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output92 (.A(net915),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output93 (.A(net916),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(clknet_1_1__leaf_net917),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net952),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output96 (.A(net919),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(clknet_1_1__leaf_net920),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(clknet_1_0__leaf_net921),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net922),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output100 (.A(net923),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_2 output101 (.A(clknet_1_1__leaf_net924),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output102 (.A(net925),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net926),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output104 (.A(net927),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output105 (.A(net928),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output106 (.A(net929),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output107 (.A(net930),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output108 (.A(net931),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output109 (.A(net932),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(clknet_1_0__leaf_net933),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net934),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output112 (.A(net935),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net936),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(clknet_1_1__leaf_net937),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net938),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(clknet_1_0__leaf_net939),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(clknet_1_1__leaf_net940),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net429),
    .X(net941));
 sky130_fd_sc_hd__buf_1 wire119 (.A(net219),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net430),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_1 max_cap121 (.A(net430),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net235),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net217),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(net217),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(net896),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_2 max_cap126 (.A(net113),
    .X(net949));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net210),
    .X(net950));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net918),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_8 fanout129 (.A(net918),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_1 max_cap130 (.A(net361),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_1 max_cap131 (.A(net141),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_1 max_cap132 (.A(net137),
    .X(net955));
 sky130_fd_sc_hd__buf_1 max_cap133 (.A(net40),
    .X(net956));
 sky130_fd_sc_hd__buf_4 max_cap134 (.A(net30),
    .X(net957));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net909),
    .X(net958));
 sky130_fd_sc_hd__buf_1 wire136 (.A(net20),
    .X(net959));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net15),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net546),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_1 max_cap140 (.A(net1005),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_2 max_cap141 (.A(net248),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_4 fanout142 (.A(net441),
    .X(net965));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(net350),
    .X(net966));
 sky130_fd_sc_hd__buf_8 fanout144 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__buf_12 fanout145 (.A(net345),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net970),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net117),
    .X(net970));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net822),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net6),
    .X(net972));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net93),
    .X(net973));
 sky130_fd_sc_hd__buf_2 max_cap151 (.A(net88),
    .X(net974));
 sky130_fd_sc_hd__inv_1 c537_1 (.A(net746),
    .Y(net975));
 sky130_fd_sc_hd__inv_1 net899_2 (.A(net746),
    .Y(net976));
 sky130_fd_sc_hd__inv_1 net899_3 (.A(net746),
    .Y(net977));
 sky130_fd_sc_hd__clkinv_2 c501_5 (.A(clknet_1_1__leaf_net748),
    .Y(net979));
 sky130_fd_sc_hd__clkinv_2 c501_6 (.A(clknet_1_0__leaf_net748),
    .Y(net980));
 sky130_fd_sc_hd__clkinv_2 c501_7 (.A(clknet_1_0__leaf_net748),
    .Y(net981));
 sky130_fd_sc_hd__clkinv_2 c501_8 (.A(clknet_1_0__leaf_net748),
    .Y(net982));
 sky130_fd_sc_hd__clkinv_2 c501_9 (.A(clknet_1_0__leaf_net748),
    .Y(net983));
 sky130_fd_sc_hd__clkinv_2 c501_10 (.A(clknet_1_0__leaf_net748),
    .Y(net984));
 sky130_fd_sc_hd__clkinv_2 c501_11 (.A(clknet_1_0__leaf_net748),
    .Y(net985));
 sky130_fd_sc_hd__clkinv_2 c501_12 (.A(clknet_1_1__leaf_net748),
    .Y(net986));
 sky130_fd_sc_hd__inv_2 c201_14 (.A(clknet_1_1__leaf_net776),
    .Y(net988));
 sky130_fd_sc_hd__inv_2 c201_15 (.A(clknet_1_1__leaf_net776),
    .Y(net989));
 sky130_fd_sc_hd__inv_2 c201_16 (.A(clknet_1_1__leaf_net776),
    .Y(net990));
 sky130_fd_sc_hd__inv_2 c201_17 (.A(clknet_1_1__leaf_net776),
    .Y(net991));
 sky130_fd_sc_hd__inv_2 c201_18 (.A(clknet_1_0__leaf_net776),
    .Y(net992));
 sky130_fd_sc_hd__inv_2 c201_19 (.A(clknet_1_0__leaf_net776),
    .Y(net993));
 sky130_fd_sc_hd__inv_2 c201_20 (.A(clknet_1_0__leaf_net776),
    .Y(net994));
 sky130_fd_sc_hd__clkinv_1 c301_22 (.A(clknet_1_0__leaf_net776),
    .Y(net996));
 sky130_fd_sc_hd__clkinv_1 c301_23 (.A(clknet_1_0__leaf_net776),
    .Y(net997));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net814 (.A(net814),
    .X(clknet_0_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net814 (.A(clknet_0_net814),
    .X(clknet_1_0__leaf_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net814 (.A(clknet_0_net814),
    .X(clknet_1_1__leaf_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net599 (.A(net599),
    .X(clknet_0_net599));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net599 (.A(clknet_0_net599),
    .X(clknet_1_0__leaf_net599));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net599 (.A(clknet_0_net599),
    .X(clknet_1_1__leaf_net599));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net598 (.A(net598),
    .X(clknet_0_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_0__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_1__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net813 (.A(net813),
    .X(clknet_0_net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net813 (.A(clknet_0_net813),
    .X(clknet_1_0__leaf_net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net813 (.A(clknet_0_net813),
    .X(clknet_1_1__leaf_net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net812 (.A(net812),
    .X(clknet_0_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net812 (.A(clknet_0_net812),
    .X(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net812 (.A(clknet_0_net812),
    .X(clknet_1_1__leaf_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net940 (.A(net940),
    .X(clknet_0_net940));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net940 (.A(net1032),
    .X(clknet_1_0__leaf_net940));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net940 (.A(clknet_0_net940),
    .X(clknet_1_1__leaf_net940));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net638 (.A(net638),
    .X(clknet_0_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net638 (.A(clknet_0_net638),
    .X(clknet_1_0__leaf_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net638 (.A(clknet_0_net638),
    .X(clknet_1_1__leaf_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net643 (.A(net643),
    .X(clknet_0_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_0__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_1__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net904 (.A(net904),
    .X(clknet_0_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net795 (.A(net795),
    .X(clknet_0_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net795 (.A(clknet_0_net795),
    .X(clknet_1_0__leaf_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net795 (.A(clknet_0_net795),
    .X(clknet_1_1__leaf_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net901 (.A(net901),
    .X(clknet_0_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net182 (.A(net182),
    .X(clknet_0_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net776 (.A(net776),
    .X(clknet_0_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net776 (.A(clknet_0_net776),
    .X(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net776 (.A(clknet_0_net776),
    .X(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net135 (.A(net135),
    .X(clknet_0_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net135 (.A(clknet_0_net135),
    .X(clknet_1_0__leaf_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net135 (.A(clknet_0_net135),
    .X(clknet_1_1__leaf_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net894 (.A(net894),
    .X(clknet_0_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net933 (.A(net933),
    .X(clknet_0_net933));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net933 (.A(clknet_0_net933),
    .X(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net933 (.A(clknet_0_net933),
    .X(clknet_1_1__leaf_net933));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net292 (.A(net292),
    .X(clknet_0_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_0__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_1__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net286 (.A(net286),
    .X(clknet_0_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_0__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_1__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net748 (.A(net748),
    .X(clknet_0_net748));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net748 (.A(clknet_0_net748),
    .X(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net748 (.A(clknet_0_net748),
    .X(clknet_1_1__leaf_net748));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net414 (.A(net414),
    .X(clknet_0_net414));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net414 (.A(clknet_0_net414),
    .X(clknet_1_0__leaf_net414));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net414 (.A(clknet_0_net414),
    .X(clknet_1_1__leaf_net414));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net423 (.A(net423),
    .X(clknet_0_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_0__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_1__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net905 (.A(net905),
    .X(clknet_0_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_0__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_1__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net937 (.A(net937),
    .X(clknet_0_net937));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net937 (.A(clknet_0_net937),
    .X(clknet_1_0__leaf_net937));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net937 (.A(clknet_0_net937),
    .X(clknet_1_1__leaf_net937));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net777 (.A(net777),
    .X(clknet_0_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_0__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_1__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net291 (.A(net291),
    .X(clknet_0_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net747 (.A(net747),
    .X(clknet_0_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_0__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_1__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net407 (.A(net407),
    .X(clknet_0_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net394 (.A(net394),
    .X(clknet_0_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_0__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_1__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net276 (.A(net276),
    .X(clknet_0_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_0__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_1__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net148 (.A(net148),
    .X(clknet_0_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net148 (.A(clknet_0_net148),
    .X(clknet_1_0__leaf_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net148 (.A(clknet_0_net148),
    .X(clknet_1_1__leaf_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net145 (.A(net145),
    .X(clknet_0_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_1__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net146 (.A(net146),
    .X(clknet_0_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net146 (.A(clknet_0_net146),
    .X(clknet_1_0__leaf_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net146 (.A(clknet_0_net146),
    .X(clknet_1_1__leaf_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net140 (.A(net140),
    .X(clknet_0_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_0__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net153 (.A(net153),
    .X(clknet_0_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net169 (.A(net169),
    .X(clknet_0_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net921 (.A(net921),
    .X(clknet_0_net921));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net921 (.A(clknet_0_net921),
    .X(clknet_1_0__leaf_net921));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net921 (.A(clknet_0_net921),
    .X(clknet_1_1__leaf_net921));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net143 (.A(net143),
    .X(clknet_0_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_0__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_1__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net395 (.A(net395),
    .X(clknet_0_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net395 (.A(clknet_0_net395),
    .X(clknet_1_0__leaf_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net395 (.A(clknet_0_net395),
    .X(clknet_1_1__leaf_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net939 (.A(net939),
    .X(clknet_0_net939));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net939 (.A(clknet_0_net939),
    .X(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net939 (.A(clknet_0_net939),
    .X(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net152 (.A(net152),
    .X(clknet_0_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net152 (.A(clknet_0_net152),
    .X(clknet_1_0__leaf_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net152 (.A(clknet_0_net152),
    .X(clknet_1_1__leaf_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net136 (.A(net136),
    .X(clknet_0_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net136 (.A(clknet_0_net136),
    .X(clknet_1_0__leaf_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net136 (.A(clknet_0_net136),
    .X(clknet_1_1__leaf_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net406 (.A(net406),
    .X(clknet_0_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_0__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_1__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net516 (.A(net516),
    .X(clknet_0_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_0__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_1__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net910 (.A(net910),
    .X(clknet_0_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_0__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_1__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net920 (.A(net920),
    .X(clknet_0_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net920 (.A(clknet_0_net920),
    .X(clknet_1_0__leaf_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net920 (.A(clknet_0_net920),
    .X(clknet_1_1__leaf_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net306 (.A(net306),
    .X(clknet_0_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_0__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_1__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net425 (.A(net425),
    .X(clknet_0_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_0__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_1__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net794 (.A(net794),
    .X(clknet_0_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net564 (.A(net564),
    .X(clknet_0_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_0__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_1__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net584 (.A(net584),
    .X(clknet_0_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_0__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net575 (.A(net575),
    .X(clknet_0_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_1__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net570 (.A(net570),
    .X(clknet_0_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net570 (.A(clknet_0_net570),
    .X(clknet_1_0__leaf_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net570 (.A(clknet_0_net570),
    .X(clknet_1_1__leaf_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net387 (.A(net387),
    .X(clknet_0_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_0__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_1__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net371 (.A(net371),
    .X(clknet_0_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_0__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_1__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net366 (.A(net366),
    .X(clknet_0_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_0__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net527 (.A(net527),
    .X(clknet_0_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_0__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_1__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net917 (.A(net917),
    .X(clknet_0_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net917 (.A(clknet_0_net917),
    .X(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net917 (.A(clknet_0_net917),
    .X(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net382 (.A(net382),
    .X(clknet_0_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_1__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net363 (.A(net363),
    .X(clknet_0_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net460 (.A(net460),
    .X(clknet_0_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_0__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_1__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net452 (.A(net452),
    .X(clknet_0_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_0__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_1__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net439 (.A(net439),
    .X(clknet_0_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_0__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_1__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net552 (.A(net552),
    .X(clknet_0_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net552 (.A(clknet_0_net552),
    .X(clknet_1_0__leaf_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net552 (.A(clknet_0_net552),
    .X(clknet_1_1__leaf_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net440 (.A(net440),
    .X(clknet_0_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_0__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_1__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net478 (.A(net478),
    .X(clknet_0_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_0__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_1__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net477 (.A(net477),
    .X(clknet_0_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_0__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_1__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net472 (.A(net472),
    .X(clknet_0_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_0__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_1__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net447 (.A(net447),
    .X(clknet_0_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_0__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_1__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net442 (.A(net442),
    .X(clknet_0_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_0__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_1__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net445 (.A(net445),
    .X(clknet_0_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_0__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_1__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net438 (.A(net438),
    .X(clknet_0_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_0__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_1__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net899 (.A(net899),
    .X(clknet_0_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net899 (.A(clknet_0_net899),
    .X(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net899 (.A(clknet_0_net899),
    .X(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net379 (.A(net379),
    .X(clknet_0_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_1__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net373 (.A(net373),
    .X(clknet_0_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_1__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net254 (.A(net254),
    .X(clknet_0_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_0__leaf_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_1__leaf_net254));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net78),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net78),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net227),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net436),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(net773),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net998),
    .X(net999));
 sky130_fd_sc_hd__buf_8 rebuffer7 (.A(net1002),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1000),
    .X(net1001));
 sky130_fd_sc_hd__buf_6 rebuffer9 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__buf_6 rebuffer10 (.A(net773),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net911),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net328),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net774),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net780),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net466),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net751),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net922),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net512),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net906),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net752),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net376),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net800),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net735),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net699),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net130),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net367),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net791),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(net141),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_1 wire2 (.A(net509),
    .X(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_C (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_Y (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_C (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_C (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_C1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_S0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_C1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_Q_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_C1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_Q (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_D1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_C_N (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_Y (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_D1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_SCE (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_C_N (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_SCD (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_Y (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_Q (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_Y (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_D_N (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_D_N (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B_N (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_Y (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_Y (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B_N (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_SCD (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Y (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_C (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_C (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_C1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_C_N (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_D1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_S1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_SCE (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_C_N (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Y (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A3 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_S1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A0 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S0 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A3 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_X (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_D1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_C (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_Q (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_Y (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_D (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_S1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_S0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_SCE (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q_N (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_C1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_SCD (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_C (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_Y (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_S1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_C (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_D_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_Y (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap134_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A_N (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_Y (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_C_N (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_D1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_B (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_B (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Y (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_S1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_SCE (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_Q_N (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_Q (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Q_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Q (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_C1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Y (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SCD (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_SCD (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_X (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_C_N (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_SCD (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_SET_B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A_N (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B_N (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_C (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_D (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_Y (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_SCD (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_SET_B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_C_N (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_C (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_D_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_C1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_C1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_Y (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B_N (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_X (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_Q_N (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_A2 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A2 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_SCD (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_C_N (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_Y (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net395_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_X (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SET_B (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_Q_N (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_Q (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_C1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_X (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_X (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_S0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_D1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_C (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_Y (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_SCE (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SCD (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_Y (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge904_D (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_X (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge906_D (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_Y (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_B (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_C1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_SET_B (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_C_N (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_C1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_Q (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_Q (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_Q (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge905_D (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_X (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_D_N (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_D (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_Y (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_Q_N (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_Q (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_D_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SCE (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_D_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_C_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_B1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_X (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_X (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_X (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A0 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S0 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_X (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_C1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_C1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_X (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_C1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_Q (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge915_RESET_B (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_Y (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_Y (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_B (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_X (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_C_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_C_N (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_C (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_D_N (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_C (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_C (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B_N (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_C_N (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_D (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Y (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B_N (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_C (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A3 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_S1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_C1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_Q (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_C (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_D1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_B_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_C_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_SCD (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold22_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q_N (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_D_N (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_Q (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_Q (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge893_Q (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge895_Q_N (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCE (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge899_Q (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_C1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_C_N (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge901_Q (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_C_N (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_C_N (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_B_N (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold19_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge904_Q (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_B1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge905_Q (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_D_N (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_D1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net776_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge907_GCLK (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_Q (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SET_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_C (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge913_Q (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_B1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge915_Q (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_B1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_D_N (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_B (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_D1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_C_N (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold33_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_Q (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q_N (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_D_N (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B_N (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_D1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_Y (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_C_N (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_Q (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_C1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SET_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_Q (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_D_N (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_Y (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_SCE (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_Y (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_Y (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SET_B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_Y (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_D (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_SCE (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_D1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C_N (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Y (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_DE (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A_N (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_D_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_C_N (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_D_N (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_D_N (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A_N (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_C (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A_N (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B_N (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_SCD (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_D1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_C1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B_N (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_C_N (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_C_N (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_B1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C_N (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B_N (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_C_N (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_C1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_C_N (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A2 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_B1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_C1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_C_N (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_SCD (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_C (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_C (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_C_N (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_D_N (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_C1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_C1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S0 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_B1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A_N (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A_N (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_C1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_D_N (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_B1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_C_N (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_Q (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge906_Q (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge905_Q_N (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_C1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_RESET_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net894_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_Q (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_C (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_Y (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_S0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_C_N (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_Y (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A_N (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_Y (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net899_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_D_N (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_D1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_Q (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_C_N (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold25_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_Q (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_C1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_D_N (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold17_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge892_Q (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_D1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_C_N (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_Q (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_Q (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge914_Q (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_D_N (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_C1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_B (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_B (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_C1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_Q (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_SCE (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_C_N (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_B (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_C_N (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_C (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_C1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_Y (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_B1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_Y (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_Q (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_C (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_Q (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_Q (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net939_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_D (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_DE (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_D (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_C1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SCE (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_B1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_B1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_C1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_C1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_C (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_C (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_D1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_D_N (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_C1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_D_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_C_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_D1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_D1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C_N (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_C_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_C_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_D_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_D1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_D1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_C_N (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_D_N (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SCE (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_B1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_C (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_C_N (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_C (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_D1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_B1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_C_N (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_D_N (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_C_N (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_D_N (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_C (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_C_N (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_C (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_C1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_D1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_C1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_C (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B_N (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_B (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B_N (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_D1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_C (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_C1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_SCE (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_C1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_C1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_C (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_SCE (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_D (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_C_N (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_C_N (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_SCE (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_D_N (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_SCE (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_C1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_B (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_D_N (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_C (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge901_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge894_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge899_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge903_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge914_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge913_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge908_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge892_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge893_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge898_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge906_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge911_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge916_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(clknet_1_1__leaf_net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net940_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net776_A (.DIODE(clknet_0_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net776_A (.DIODE(clknet_0_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net776_X (.DIODE(clknet_0_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_C (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_D1 (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_D1 (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_18_A (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_19_A (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_20_A (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_21_A (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_22_A (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_23_A (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net776_X (.DIODE(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_C1 (.DIODE(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_13_A (.DIODE(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_14_A (.DIODE(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_15_A (.DIODE(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_16_A (.DIODE(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_17_A (.DIODE(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net776_X (.DIODE(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net894_A (.DIODE(clknet_0_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net894_A (.DIODE(clknet_0_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net894_X (.DIODE(clknet_0_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S0 (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_D1 (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A2 (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A2 (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net894_X (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_C1 (.DIODE(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_SET_B (.DIODE(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net894_X (.DIODE(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_C_N (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_C1 (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A2 (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A2 (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net933_X (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_6_A (.DIODE(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_7_A (.DIODE(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_8_A (.DIODE(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_9_A (.DIODE(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_10_A (.DIODE(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_11_A (.DIODE(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net748_X (.DIODE(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_C (.DIODE(clknet_1_1__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A (.DIODE(clknet_1_1__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_4_A (.DIODE(clknet_1_1__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_5_A (.DIODE(clknet_1_1__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_12_A (.DIODE(clknet_1_1__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net748_X (.DIODE(clknet_1_1__leaf_net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_SCD (.DIODE(clknet_1_0__leaf_net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A2 (.DIODE(clknet_1_0__leaf_net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(clknet_1_0__leaf_net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net921_X (.DIODE(clknet_1_0__leaf_net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_B1 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_D1 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A3 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_SCD (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A3 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_C_N (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net939_X (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_SET_B (.DIODE(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_SCD (.DIODE(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SCD (.DIODE(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net939_X (.DIODE(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_D1 (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_C_N (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_D1 (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_D_N (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SCE (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net794_X (.DIODE(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_D1 (.DIODE(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_D_N (.DIODE(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_D_N (.DIODE(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_D_N (.DIODE(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_D1 (.DIODE(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net794_X (.DIODE(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_B1 (.DIODE(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net584_X (.DIODE(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_RESET_B (.DIODE(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net365_X (.DIODE(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net899_A (.DIODE(clknet_0_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net899_A (.DIODE(clknet_0_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net899_X (.DIODE(clknet_0_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B1 (.DIODE(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B1 (.DIODE(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_D1 (.DIODE(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C1 (.DIODE(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B1 (.DIODE(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_D (.DIODE(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net899_X (.DIODE(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A3 (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A2 (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net899_X (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(clknet_1_0__leaf_net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A1 (.DIODE(clknet_1_0__leaf_net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net254_X (.DIODE(clknet_1_0__leaf_net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_C1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_X (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net951));
 sky130_fd_sc_hd__nor2b_1 clone1 (.A(net64),
    .B_N(net824),
    .Y(net1006));
 sky130_fd_sc_hd__or3_1 clone2 (.A(net343),
    .B(net65),
    .C(net967),
    .X(net1007));
 sky130_fd_sc_hd__or2b_1 clone3 (.A(net67),
    .B_N(net825),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net69),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_1 clone12 (.A(net345),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net191),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1028),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net1028),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_1 clone16 (.A(clknet_0_net940),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(clknet_0_net940),
    .X(net1032));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
