module netlist_1 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input in52,
	input in53,
	input in54,
	input in55,
	input in56,
	input in57,
	input in58,
	input in59,
	input in60,
	input in61,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51,
	output out52,
	output out53,
	output out54,
	output out55,
	output out56,
	output out57,
	output out58,
	output out59,
	output out60,
	output out61
);


wire clk;
wire net766;
wire net765;
wire net764;
wire net763;
wire net762;
wire net759;
wire net755;
wire net754;
wire net753;
wire net752;
wire net751;
wire net750;
wire net748;
wire net747;
wire net745;
wire net744;
wire net743;
wire net741;
wire net740;
wire net739;
wire net738;
wire net735;
wire net732;
wire net731;
wire net730;
wire net729;
wire net728;
wire net726;
wire net725;
wire net724;
wire out15;
wire net722;
wire out18;
wire net720;
wire net719;
wire net717;
wire net716;
wire net715;
wire net714;
wire net712;
wire net711;
wire net708;
wire net706;
wire net705;
wire net704;
wire net703;
wire out32;
wire net701;
wire net699;
wire net698;
wire net697;
wire net696;
wire net695;
wire net694;
wire net693;
wire net692;
wire net690;
wire out8;
wire net687;
wire net686;
wire out24;
wire net685;
wire net684;
wire net683;
wire out57;
wire net503;
wire net679;
wire net671;
wire net669;
wire net668;
wire net370;
wire net667;
wire net664;
wire net659;
wire in6;
wire net656;
wire net652;
wire net622;
wire net651;
wire net304;
wire net645;
wire net641;
wire net637;
wire net632;
wire net665;
wire net631;
wire net629;
wire net74;
wire net628;
wire net3;
wire net627;
wire net447;
wire net626;
wire net624;
wire net506;
wire net623;
wire net620;
wire in49;
wire net619;
wire net46;
wire net615;
wire net100;
wire net347;
wire net288;
wire net614;
wire net165;
wire net613;
wire net20;
wire net612;
wire net638;
wire net428;
wire net610;
wire out25;
wire net608;
wire net1;
wire net424;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire net596;
wire net592;
wire net588;
wire net587;
wire in4;
wire net583;
wire net707;
wire net582;
wire net158;
wire net584;
wire net581;
wire net336;
wire net579;
wire net577;
wire net576;
wire net209;
wire net569;
wire in41;
wire net567;
wire in30;
wire net566;
wire net565;
wire net39;
wire net562;
wire net559;
wire net556;
wire net647;
wire net555;
wire net159;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire in55;
wire net550;
wire net710;
wire net544;
wire net539;
wire net534;
wire net532;
wire net271;
wire net530;
wire net617;
wire net306;
wire net537;
wire net369;
wire net528;
wire net525;
wire net523;
wire net520;
wire net519;
wire net516;
wire net672;
wire net514;
wire net18;
wire out34;
wire net512;
wire net78;
wire net508;
wire net721;
wire net504;
wire net224;
wire net573;
wire net499;
wire net674;
wire net496;
wire net495;
wire net494;
wire net179;
wire in39;
wire net453;
wire net493;
wire net472;
wire net492;
wire net479;
wire net491;
wire net295;
wire net490;
wire net489;
wire net487;
wire net486;
wire out1;
wire net478;
wire net474;
wire net473;
wire net468;
wire net540;
wire net202;
wire net465;
wire out7;
wire net462;
wire net469;
wire net471;
wire net461;
wire net546;
wire net749;
wire net460;
wire net454;
wire net648;
wire net452;
wire net449;
wire net448;
wire net498;
wire net700;
wire net446;
wire net680;
wire net691;
wire net88;
wire net444;
wire in59;
wire net110;
wire net442;
wire net441;
wire net609;
wire net440;
wire out11;
wire net128;
wire net439;
wire net147;
wire out21;
wire net438;
wire net433;
wire net432;
wire out41;
wire net419;
wire net431;
wire net430;
wire net618;
wire net429;
wire net427;
wire net426;
wire net673;
wire net425;
wire net423;
wire net183;
wire net531;
wire net421;
wire net52;
wire net170;
wire net420;
wire net450;
wire net418;
wire net415;
wire net414;
wire net276;
wire net413;
wire net252;
wire net330;
wire net412;
wire net411;
wire net517;
wire net677;
wire net410;
wire net409;
wire net407;
wire net662;
wire net405;
wire net607;
wire net526;
wire net404;
wire net29;
wire net403;
wire net383;
wire net663;
wire net402;
wire net106;
wire net572;
wire net401;
wire net399;
wire net398;
wire net476;
wire net396;
wire net391;
wire net443;
wire net557;
wire net345;
wire net527;
wire net488;
wire net390;
wire out5;
wire net646;
wire net389;
wire net513;
wire out14;
wire net501;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net184;
wire net131;
wire net380;
wire net379;
wire net260;
wire net616;
wire net378;
wire net543;
wire net38;
wire net377;
wire net376;
wire net625;
wire net373;
wire net598;
wire net374;
wire out20;
wire net676;
wire net372;
wire net371;
wire net368;
wire net367;
wire net366;
wire net365;
wire net364;
wire net363;
wire net360;
wire net397;
wire net357;
wire net356;
wire net510;
wire net355;
wire out6;
wire net590;
wire net507;
wire net351;
wire net746;
wire net350;
wire net547;
wire net511;
wire net451;
wire net13;
wire net343;
wire net89;
wire net666;
wire net340;
wire net339;
wire net337;
wire net458;
wire net538;
wire net244;
wire net334;
wire net333;
wire net332;
wire net331;
wire net328;
wire net327;
wire net119;
wire net325;
wire net324;
wire net321;
wire net406;
wire out19;
wire net535;
wire net320;
wire net542;
wire net139;
wire net318;
wire out31;
wire net316;
wire out9;
wire net335;
wire net315;
wire net313;
wire net505;
wire net199;
wire out27;
wire net294;
wire net319;
wire net312;
wire net742;
wire net308;
wire net352;
wire net307;
wire net305;
wire net291;
wire net303;
wire net417;
wire net302;
wire net301;
wire net298;
wire net459;
wire net463;
wire net0;
wire net297;
wire net296;
wire in24;
wire net358;
wire net127;
wire net293;
wire net292;
wire net500;
wire net445;
wire net230;
wire out22;
wire net201;
wire net422;
wire net289;
wire net595;
wire net384;
wire net482;
wire in25;
wire in8;
wire net30;
wire out36;
wire net589;
wire net278;
wire net761;
wire net274;
wire net643;
wire net273;
wire net142;
wire out10;
wire net272;
wire net757;
wire in56;
wire net134;
wire out48;
wire net114;
wire net270;
wire in17;
wire net267;
wire net644;
wire net266;
wire net408;
wire net475;
wire net280;
wire net102;
wire net151;
wire net275;
wire net264;
wire net657;
wire net591;
wire net196;
wire net262;
wire net217;
wire net261;
wire net21;
wire net257;
wire net689;
wire net44;
wire net117;
wire net62;
wire net109;
wire net254;
wire net203;
wire net253;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire in26;
wire net661;
wire net194;
wire net241;
wire net416;
wire net41;
wire net104;
wire net8;
wire out33;
wire in29;
wire net240;
wire net238;
wire net234;
wire net232;
wire out12;
wire net226;
wire net568;
wire net375;
wire net223;
wire net524;
wire net575;
wire net382;
wire net548;
wire net259;
wire net222;
wire net31;
wire net219;
wire net578;
wire net210;
wire net326;
wire net213;
wire net208;
wire out16;
wire net188;
wire net207;
wire net649;
wire net205;
wire net521;
wire net353;
wire net678;
wire net633;
wire net122;
wire net197;
wire net483;
wire net193;
wire net192;
wire net737;
wire net190;
wire net630;
wire in20;
wire net189;
wire net246;
wire net186;
wire net152;
wire net126;
wire net113;
wire net284;
wire net655;
wire net563;
wire net464;
wire net549;
wire net182;
wire net310;
wire net180;
wire out40;
wire net258;
wire out23;
wire net176;
wire net580;
wire net133;
wire net175;
wire net80;
wire net173;
wire out52;
wire net195;
wire net395;
wire net172;
wire net342;
wire net17;
wire net437;
wire out44;
wire in37;
wire net518;
wire net381;
wire net218;
wire net300;
wire net169;
wire net485;
wire net344;
wire net168;
wire net153;
wire net286;
wire net167;
wire net509;
wire net58;
wire net221;
wire net166;
wire net269;
wire out60;
wire net497;
wire net161;
wire net285;
wire net160;
wire net636;
wire net311;
wire net767;
wire net111;
wire net124;
wire net242;
wire net290;
wire net227;
wire out47;
wire net150;
wire net149;
wire net148;
wire net178;
wire net239;
wire net144;
wire net322;
wire net688;
wire net299;
wire net758;
wire net143;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net561;
wire net137;
wire net136;
wire net456;
wire net135;
wire net255;
wire net157;
wire net177;
wire net349;
wire out51;
wire net250;
wire net225;
wire net132;
wire out49;
wire out61;
wire net130;
wire net481;
wire net120;
wire net200;
wire net204;
wire out17;
wire out0;
wire net164;
wire net642;
wire net268;
wire in7;
wire net756;
wire net400;
wire net82;
wire net2;
wire net123;
wire net282;
wire net71;
wire net229;
wire in43;
wire net108;
wire net107;
wire net660;
wire net359;
wire out28;
wire in12;
wire net103;
wire out26;
wire net99;
wire net348;
wire net341;
wire in52;
wire net96;
wire net466;
wire net118;
wire net94;
wire net90;
wire net174;
wire net277;
wire net639;
wire net81;
wire in10;
wire net156;
wire net361;
wire net115;
wire net670;
wire in18;
wire net27;
wire net34;
wire net585;
wire net79;
wire net231;
wire net329;
wire net212;
wire net653;
wire in5;
wire net14;
wire net77;
wire net600;
wire net236;
wire net76;
wire in42;
wire net354;
wire in38;
wire net736;
wire net198;
wire net467;
wire net101;
wire net9;
wire net75;
wire out50;
wire net457;
wire net42;
wire net91;
wire out4;
wire net571;
wire net73;
wire net116;
wire net69;
wire net67;
wire net98;
wire net522;
wire net436;
wire net541;
wire net323;
wire net15;
wire net279;
wire net64;
wire net63;
wire net681;
wire net61;
wire net60;
wire net564;
wire net154;
wire net84;
wire net237;
wire net682;
wire in46;
wire net85;
wire net72;
wire net392;
wire out37;
wire net97;
wire net434;
wire net621;
wire net162;
wire out3;
wire net59;
wire net248;
wire net477;
wire net228;
wire net675;
wire net56;
wire out53;
wire net55;
wire net214;
wire net53;
wire in48;
wire out56;
wire out38;
wire net640;
wire net50;
wire net597;
wire out55;
wire net185;
wire net155;
wire net338;
wire net599;
wire net112;
wire net650;
wire net560;
wire net45;
wire net502;
wire net235;
wire net49;
wire net594;
wire in50;
wire net215;
wire net484;
wire net346;
wire net4;
wire net43;
wire net233;
wire net33;
wire net187;
wire in13;
wire net586;
wire net533;
wire net32;
wire net125;
wire net19;
wire in15;
wire net727;
wire net163;
wire in19;
wire net702;
wire net70;
wire net48;
wire net28;
wire net92;
wire net713;
wire net25;
wire net570;
wire out2;
wire in0;
wire out59;
wire net709;
wire net24;
wire net470;
wire in33;
wire net40;
wire in60;
wire net435;
wire net760;
wire net23;
wire net26;
wire net16;
wire in31;
wire net129;
wire net65;
wire in32;
wire net601;
wire out35;
wire net558;
wire in1;
wire net265;
wire net22;
wire net263;
wire net6;
wire net5;
wire net206;
wire in58;
wire in61;
wire net733;
wire net171;
wire in23;
wire in57;
wire net281;
wire net54;
wire in54;
wire in53;
wire net138;
wire net145;
wire net211;
wire in35;
wire in34;
wire net593;
wire in45;
wire net393;
wire net256;
wire net87;
wire net181;
wire net7;
wire out54;
wire net574;
wire net216;
wire net455;
wire in28;
wire in44;
wire net47;
wire net12;
wire in27;
wire in9;
wire net654;
wire net723;
wire net611;
wire net515;
wire net362;
wire in16;
wire out46;
wire net191;
wire net35;
wire net309;
wire net220;
wire in22;
wire net68;
wire in14;
wire net529;
wire in21;
wire net57;
wire net480;
wire net86;
wire net317;
wire in51;
wire net93;
wire in47;
wire in2;
wire net718;
wire net658;
wire net105;
wire out13;
wire in11;
wire net51;
wire out30;
wire in36;
wire net536;
wire net37;
wire net36;
wire net95;
wire net121;
wire net146;
wire net734;
wire net251;
wire net768;
wire net11;
wire net394;
wire net314;
wire in3;
wire out58;
sky130_fd_sc_hd__mux4_4 c62(
.A0(in44),
.A1(in55),
.A2(in53),
.A3(in52),
.S0(in49),
.S1(in58),
.X(net0)
);

sky130_fd_sc_hd__mux4_4 c63(
.A0(in50),
.A1(in44),
.A2(in53),
.A3(in49),
.S0(in38),
.S1(in48),
.X(net1)
);

sky130_fd_sc_hd__mux4_1 c64(
.A0(in32),
.A1(in14),
.A2(in38),
.A3(in53),
.S0(in57),
.S1(in52),
.X(net2)
);

sky130_fd_sc_hd__o211a_1 c65(
.A1(in35),
.A2(in39),
.B1(in32),
.C1(in26),
.X(net3)
);

sky130_fd_sc_hd__nor2_2 c66(
.A(net3),
.B(in25),
.Y(net4)
);

sky130_fd_sc_hd__or2_4 c67(
.A(net2),
.B(in38),
.X(net5)
);

sky130_fd_sc_hd__and2b_2 c68(
.A_N(in51),
.B(in9),
.X(net6)
);

sky130_fd_sc_hd__or2b_1 c69(
.A(net4),
.B_N(net6),
.X(net7)
);

sky130_fd_sc_hd__or2_1 c70(
.A(in44),
.B(net4),
.X(out12)
);

sky130_fd_sc_hd__or2b_4 c71(
.A(in22),
.B_N(out12),
.X(net8)
);

sky130_fd_sc_hd__nand2_1 c72(
.A(net6),
.B(in22),
.Y(net9)
);

sky130_fd_sc_hd__nand2b_2 c73(
.A_N(net1),
.B(in25),
.Y(net10)
);

sky130_fd_sc_hd__nor2b_1 c74(
.A(net5),
.B_N(net6),
.Y(net11)
);

sky130_fd_sc_hd__nor3_1 c75(
.A(out12),
.B(in44),
.C(net11),
.Y(net12)
);

sky130_fd_sc_hd__and2b_2 c76(
.A_N(net11),
.B(net12),
.X(net13)
);

sky130_fd_sc_hd__and2_4 c77(
.A(in18),
.B(in45),
.X(net14)
);

sky130_fd_sc_hd__or2b_4 c78(
.A(net13),
.B_N(out12),
.X(out35)
);

sky130_fd_sc_hd__nand3_2 c79(
.A(in56),
.B(net5),
.C(net11),
.Y(out53)
);

sky130_fd_sc_hd__nand2_4 c80(
.A(net10),
.B(net14),
.Y(net15)
);

sky130_fd_sc_hd__or2_2 c81(
.A(in43),
.B(net11),
.X(net16)
);

sky130_fd_sc_hd__mux4_1 c82(
.A0(net15),
.A1(net11),
.A2(in16),
.A3(net7),
.S0(net4),
.S1(out12),
.X(net17)
);

sky130_fd_sc_hd__mux4_4 c83(
.A0(net14),
.A1(net15),
.A2(net13),
.A3(in43),
.S0(out35),
.S1(net9),
.X(net18)
);

sky130_fd_sc_hd__nor2b_4 c84(
.A(net16),
.B_N(net17),
.Y(net19)
);

sky130_fd_sc_hd__and3_2 c85(
.A(net18),
.B(net16),
.C(net15),
.X(net20)
);

sky130_fd_sc_hd__o221a_2 c86(
.A1(net20),
.A2(net16),
.B1(net17),
.B2(out12),
.C1(out35),
.X(net21)
);

sky130_fd_sc_hd__or3b_2 c87(
.A(net8),
.B(net12),
.C_N(net21),
.X(net22)
);

sky130_fd_sc_hd__nand2b_2 c88(
.A_N(net5),
.B(net18),
.Y(net23)
);

sky130_fd_sc_hd__nand2b_4 c89(
.A_N(net7),
.B(net0),
.Y(net24)
);

sky130_fd_sc_hd__or2b_2 c90(
.A(in26),
.B_N(out35),
.X(net25)
);

sky130_fd_sc_hd__and2_2 c91(
.A(net15),
.B(net8),
.X(net26)
);

sky130_fd_sc_hd__and2b_1 c92(
.A_N(in38),
.B(in48),
.X(net27)
);

sky130_fd_sc_hd__nand2b_4 c93(
.A_N(net1),
.B(net25),
.Y(net28)
);

sky130_fd_sc_hd__and2b_4 c94(
.A_N(net25),
.B(net27),
.X(net29)
);

sky130_fd_sc_hd__nand3_2 c95(
.A(net28),
.B(net24),
.C(net25),
.Y(net30)
);

sky130_fd_sc_hd__or3_4 c96(
.A(net27),
.B(net30),
.C(net29),
.X(net31)
);

sky130_fd_sc_hd__o211ai_4 c97(
.A1(net24),
.A2(net18),
.B1(net25),
.C1(in48),
.Y(net32)
);

sky130_fd_sc_hd__and3_2 c98(
.A(net23),
.B(out53),
.C(net30),
.X(net33)
);

sky130_fd_sc_hd__nand3_2 c99(
.A(net28),
.B(net27),
.C(net29),
.Y(net34)
);

sky130_fd_sc_hd__o211a_1 c100(
.A1(in20),
.A2(net32),
.B1(net30),
.C1(net7),
.X(net35)
);

sky130_fd_sc_hd__or3b_2 c101(
.A(net29),
.B(net31),
.C_N(net33),
.X(net36)
);

sky130_fd_sc_hd__and3b_1 c102(
.A_N(net31),
.B(net32),
.C(net28),
.X(net37)
);

sky130_fd_sc_hd__mux4_4 c103(
.A0(net35),
.A1(net34),
.A2(net23),
.A3(net37),
.S0(net30),
.S1(net24),
.X(net38)
);

sky130_fd_sc_hd__and3b_2 c104(
.A_N(net37),
.B(net36),
.C(net18),
.X(net39)
);

sky130_fd_sc_hd__mux4_4 c105(
.A0(net39),
.A1(net29),
.A2(net27),
.A3(net28),
.S0(in26),
.S1(net38),
.X(net40)
);

sky130_fd_sc_hd__mux4_1 c106(
.A0(in38),
.A1(net12),
.A2(net37),
.A3(net39),
.S0(net29),
.S1(net40),
.X(net41)
);

sky130_fd_sc_hd__o221a_1 c107(
.A1(net32),
.A2(net37),
.B1(net39),
.B2(net38),
.C1(net34),
.X(net42)
);

sky130_fd_sc_hd__and3_4 c108(
.A(net33),
.B(net39),
.C(net42),
.X(net43)
);

sky130_fd_sc_hd__mux4_4 c109(
.A0(net40),
.A1(net43),
.A2(net36),
.A3(net30),
.S0(net42),
.S1(net41),
.X(net44)
);

sky130_fd_sc_hd__nor2_2 c110(
.A(in19),
.B(net24),
.Y(net45)
);

sky130_fd_sc_hd__nor2_1 c111(
.A(net4),
.B(net29),
.Y(net46)
);

sky130_fd_sc_hd__nor3b_2 c112(
.A(net45),
.B(in0),
.C_N(net24),
.Y(net47)
);

sky130_fd_sc_hd__nor2b_4 c113(
.A(net16),
.B_N(net46),
.Y(net48)
);

sky130_fd_sc_hd__nand2_4 c114(
.A(net8),
.B(net24),
.Y(net49)
);

sky130_fd_sc_hd__o221a_1 c115(
.A1(net49),
.A2(net46),
.B1(net29),
.B2(net47),
.C1(net48),
.X(net50)
);

sky130_fd_sc_hd__o221ai_4 c116(
.A1(net45),
.A2(net29),
.B1(net43),
.B2(net24),
.C1(net39),
.Y(net51)
);

sky130_fd_sc_hd__and2_2 c117(
.A(net48),
.B(net4),
.X(out38)
);

sky130_fd_sc_hd__or2b_1 c118(
.A(net46),
.B_N(net51),
.X(net52)
);

sky130_fd_sc_hd__o221ai_1 c119(
.A1(net24),
.A2(net22),
.B1(out53),
.B2(out38),
.C1(net29),
.Y(net53)
);

sky130_fd_sc_hd__nor2b_2 c120(
.A(net49),
.B_N(net50),
.Y(net54)
);

sky130_fd_sc_hd__nand2b_4 c121(
.A_N(net53),
.B(net54),
.Y(net55)
);

sky130_fd_sc_hd__o211a_1 c122(
.A1(in46),
.A2(net52),
.B1(net24),
.C1(in45),
.X(net56)
);

sky130_fd_sc_hd__nand3b_1 c123(
.A_N(net55),
.B(net53),
.C(in46),
.Y(net57)
);

sky130_fd_sc_hd__mux4_2 c124(
.A0(net56),
.A1(in36),
.A2(net53),
.A3(net47),
.S0(net49),
.S1(net46),
.X(net58)
);

sky130_fd_sc_hd__o221a_4 c125(
.A1(in9),
.A2(net52),
.B1(net58),
.B2(net43),
.C1(net56),
.X(net59)
);

sky130_fd_sc_hd__o211ai_4 c126(
.A1(net54),
.A2(net57),
.B1(net45),
.C1(net55),
.Y(net60)
);

sky130_fd_sc_hd__mux4_4 c127(
.A0(net22),
.A1(net54),
.A2(net53),
.A3(net46),
.S0(net52),
.S1(net57),
.X(out3)
);

sky130_fd_sc_hd__and2_0 c128(
.A(net47),
.B(net45),
.X(out57)
);

sky130_fd_sc_hd__o221a_2 c129(
.A1(net57),
.A2(net54),
.B1(net60),
.B2(out3),
.C1(net24),
.X(out5)
);

sky130_fd_sc_hd__mux4_4 c130(
.A0(net52),
.A1(net39),
.A2(out5),
.A3(net59),
.S0(out3),
.S1(out57),
.X(net61)
);

sky130_fd_sc_hd__mux4_2 c131(
.A0(net61),
.A1(out3),
.A2(out57),
.A3(out38),
.S0(net56),
.S1(net59),
.X(net62)
);

sky130_fd_sc_hd__nor2b_4 c132(
.A(in18),
.B_N(in20),
.Y(out10)
);

sky130_fd_sc_hd__and2b_1 c133(
.A_N(out10),
.B(in13),
.X(net63)
);

sky130_fd_sc_hd__nand2_1 c134(
.A(net63),
.B(out10),
.Y(net64)
);

sky130_fd_sc_hd__nand2b_1 c135(
.A_N(in11),
.B(in16),
.Y(net65)
);

sky130_fd_sc_hd__nor2b_2 c136(
.A(in7),
.B_N(in15),
.Y(net66)
);

sky130_fd_sc_hd__nor3_4 c137(
.A(in8),
.B(in12),
.C(in4),
.Y(net67)
);

sky130_fd_sc_hd__or2_2 c138(
.A(in15),
.B(in6),
.X(net68)
);

sky130_fd_sc_hd__nand3b_4 c139(
.A_N(out10),
.B(net63),
.C(in3),
.Y(net69)
);

sky130_fd_sc_hd__nor3b_1 c140(
.A(net64),
.B(net68),
.C_N(net67),
.Y(net70)
);

sky130_fd_sc_hd__or2b_2 c141(
.A(net68),
.B_N(net64),
.X(net71)
);

sky130_fd_sc_hd__or3_4 c142(
.A(in3),
.B(net70),
.C(net63),
.X(net72)
);

sky130_fd_sc_hd__mux4_1 c143(
.A0(net63),
.A1(in11),
.A2(in21),
.A3(net72),
.S0(net68),
.S1(net70),
.X(net73)
);

sky130_fd_sc_hd__nand3_4 c144(
.A(net69),
.B(in10),
.C(net65),
.Y(net74)
);

sky130_fd_sc_hd__nor2_1 c145(
.A(net73),
.B(net67),
.Y(net75)
);

sky130_fd_sc_hd__nand3_2 c146(
.A(net71),
.B(net65),
.C(in14),
.Y(net76)
);

sky130_fd_sc_hd__nor3b_1 c147(
.A(net70),
.B(in14),
.C_N(net64),
.Y(net77)
);

sky130_fd_sc_hd__or3b_4 c148(
.A(net76),
.B(in16),
.C_N(in1),
.X(net78)
);

sky130_fd_sc_hd__o221a_2 c149(
.A1(net72),
.A2(net67),
.B1(net73),
.B2(in6),
.C1(in5),
.X(net79)
);

sky130_fd_sc_hd__or3b_1 c150(
.A(net79),
.B(out10),
.C_N(net71),
.X(net80)
);

sky130_fd_sc_hd__mux4_2 c151(
.A0(net78),
.A1(net77),
.A2(net64),
.A3(in13),
.S0(net63),
.S1(in5),
.X(net81)
);

sky130_fd_sc_hd__or3b_1 c152(
.A(in13),
.B(net80),
.C_N(net67),
.X(net82)
);

sky130_fd_sc_hd__nor3b_4 c153(
.A(net81),
.B(in21),
.C_N(net79),
.Y(net83)
);

sky130_fd_sc_hd__or2_4 c154(
.A(net72),
.B(in24),
.X(net84)
);

sky130_fd_sc_hd__or2b_2 c155(
.A(net79),
.B_N(in25),
.X(net85)
);

sky130_fd_sc_hd__and3b_1 c156(
.A_N(in41),
.B(net71),
.C(net85),
.X(net86)
);

sky130_fd_sc_hd__nand2b_1 c157(
.A_N(net71),
.B(in31),
.Y(net87)
);

sky130_fd_sc_hd__and2_4 c158(
.A(net66),
.B(in42),
.X(net88)
);

sky130_fd_sc_hd__or2b_1 c159(
.A(net82),
.B_N(in23),
.X(net89)
);

sky130_fd_sc_hd__nand2_2 c160(
.A(net87),
.B(in40),
.Y(net90)
);

sky130_fd_sc_hd__and2b_1 c161(
.A_N(net86),
.B(in34),
.X(net91)
);

sky130_fd_sc_hd__nand3b_2 c162(
.A_N(in28),
.B(net84),
.C(net91),
.Y(net92)
);

sky130_fd_sc_hd__o211ai_1 c163(
.A1(net86),
.A2(net92),
.B1(in4),
.C1(net89),
.Y(out58)
);

sky130_fd_sc_hd__o221a_2 c164(
.A1(net91),
.A2(in12),
.B1(net87),
.B2(in39),
.C1(out10),
.X(net93)
);

sky130_fd_sc_hd__nor2_4 c165(
.A(net65),
.B(in6),
.Y(net94)
);

sky130_fd_sc_hd__mux4_2 c166(
.A0(in42),
.A1(in18),
.A2(net94),
.A3(in41),
.S0(net85),
.S1(net89),
.X(net95)
);

sky130_fd_sc_hd__or3_2 c167(
.A(in40),
.B(net90),
.C(net94),
.X(net96)
);

sky130_fd_sc_hd__nand3b_1 c168(
.A_N(in26),
.B(net95),
.C(net94),
.Y(net97)
);

sky130_fd_sc_hd__or2_2 c169(
.A(net97),
.B(net94),
.X(net98)
);

sky130_fd_sc_hd__o211a_4 c170(
.A1(net96),
.A2(net89),
.B1(net97),
.C1(net94),
.X(net99)
);

sky130_fd_sc_hd__nand3b_4 c171(
.A_N(net99),
.B(net94),
.C(net89),
.Y(net100)
);

sky130_fd_sc_hd__mux4_1 c172(
.A0(net93),
.A1(net99),
.A2(net97),
.A3(net94),
.S0(in31),
.S1(in39),
.X(net101)
);

sky130_fd_sc_hd__o211a_2 c173(
.A1(net91),
.A2(net88),
.B1(net100),
.C1(net94),
.X(net102)
);

sky130_fd_sc_hd__mux4_2 c174(
.A0(in4),
.A1(net102),
.A2(net87),
.A3(net101),
.S0(net94),
.S1(net93),
.X(net103)
);

sky130_fd_sc_hd__o211ai_4 c175(
.A1(net101),
.A2(net103),
.B1(net100),
.C1(net94),
.Y(net104)
);

sky130_fd_sc_hd__or2b_2 c176(
.A(net100),
.B_N(in53),
.X(out28)
);

sky130_fd_sc_hd__or2b_2 c177(
.A(net95),
.B_N(out58),
.X(net105)
);

sky130_fd_sc_hd__and3b_2 c178(
.A_N(net83),
.B(in54),
.C(net70),
.X(net106)
);

sky130_fd_sc_hd__or2_1 c179(
.A(in1),
.B(net74),
.X(out37)
);

sky130_fd_sc_hd__and2_1 c180(
.A(in30),
.B(net91),
.X(net107)
);

sky130_fd_sc_hd__nor2_1 c181(
.A(net89),
.B(in27),
.Y(net108)
);

sky130_fd_sc_hd__and2_1 c182(
.A(in45),
.B(in52),
.X(net109)
);

sky130_fd_sc_hd__nor2_1 c183(
.A(out28),
.B(in60),
.Y(net110)
);

sky130_fd_sc_hd__nand3b_4 c184(
.A_N(in37),
.B(net83),
.C(net106),
.Y(net111)
);

sky130_fd_sc_hd__nand2b_4 c185(
.A_N(in52),
.B(net111),
.Y(net112)
);

sky130_fd_sc_hd__mux4_4 c186(
.A0(in60),
.A1(net112),
.A2(net107),
.A3(in52),
.S0(net111),
.S1(net89),
.X(net113)
);

sky130_fd_sc_hd__o211ai_4 c187(
.A1(net3),
.A2(in58),
.B1(in45),
.C1(net99),
.Y(net114)
);

sky130_fd_sc_hd__o211ai_4 c188(
.A1(net105),
.A2(out28),
.B1(net89),
.C1(net114),
.Y(net115)
);

sky130_fd_sc_hd__nand3_1 c189(
.A(net103),
.B(net100),
.C(net115),
.Y(net116)
);

sky130_fd_sc_hd__nand3_4 c190(
.A(net107),
.B(net116),
.C(net111),
.Y(net117)
);

sky130_fd_sc_hd__o211ai_1 c191(
.A1(net115),
.A2(in30),
.B1(net116),
.C1(net89),
.Y(net118)
);

sky130_fd_sc_hd__o211a_2 c192(
.A1(net108),
.A2(in1),
.B1(net117),
.C1(net66),
.X(net119)
);

sky130_fd_sc_hd__o221ai_4 c193(
.A1(net112),
.A2(net119),
.B1(net114),
.B2(out37),
.C1(in49),
.Y(net120)
);

sky130_fd_sc_hd__and2b_2 c194(
.A_N(net114),
.B(net115),
.X(net121)
);

sky130_fd_sc_hd__and3_2 c195(
.A(net115),
.B(net104),
.C(net84),
.X(net122)
);

sky130_fd_sc_hd__mux4_4 c196(
.A0(in12),
.A1(net83),
.A2(in37),
.A3(net89),
.S0(net107),
.S1(net122),
.X(net123)
);

sky130_fd_sc_hd__mux4_2 c197(
.A0(net119),
.A1(net116),
.A2(net122),
.A3(net115),
.S0(net123),
.S1(net112),
.X(net124)
);

sky130_fd_sc_hd__or3b_1 c198(
.A(net92),
.B(in45),
.C_N(net109),
.X(net125)
);

sky130_fd_sc_hd__or2_2 c199(
.A(in21),
.B(net113),
.X(net126)
);

sky130_fd_sc_hd__or2b_2 c200(
.A(net13),
.B_N(net126),
.X(net127)
);

sky130_fd_sc_hd__nand2_2 c201(
.A(in33),
.B(net124),
.Y(net128)
);

sky130_fd_sc_hd__nand2_2 c202(
.A(net123),
.B(net126),
.Y(net129)
);

sky130_fd_sc_hd__nand2b_1 c203(
.A_N(net126),
.B(net92),
.Y(net130)
);

sky130_fd_sc_hd__nor2b_2 c204(
.A(net107),
.B_N(in58),
.Y(net131)
);

sky130_fd_sc_hd__and3_4 c205(
.A(net126),
.B(net129),
.C(net10),
.X(out61)
);

sky130_fd_sc_hd__nand3b_4 c206(
.A_N(net109),
.B(net125),
.C(net127),
.Y(net132)
);

sky130_fd_sc_hd__dlygate4sd1_1 c207(
.A(net627),
.X(net133)
);

sky130_fd_sc_hd__o221a_4 c208(
.A1(net113),
.A2(net14),
.B1(net9),
.B2(out61),
.C1(net126),
.X(net134)
);

sky130_fd_sc_hd__o221ai_1 c209(
.A1(net9),
.A2(net113),
.B1(net66),
.B2(net126),
.C1(net674),
.Y(net135)
);

sky130_fd_sc_hd__nor2b_2 c210(
.A(net135),
.B_N(net127),
.Y(net136)
);

sky130_fd_sc_hd__o211a_2 c211(
.A1(net116),
.A2(in34),
.B1(in25),
.C1(net135),
.X(net137)
);

sky130_fd_sc_hd__or2b_4 c212(
.A(in25),
.B_N(net21),
.X(net138)
);

sky130_fd_sc_hd__sdfbbn_1 c213(
.D(net131),
.RESET_B(in33),
.SCD(net130),
.SCE(net13),
.SET_B(out61),
.CLK_N(clk),
.Q(net140),
.Q_N(net139)
);

sky130_fd_sc_hd__o211ai_4 c214(
.A1(net136),
.A2(net107),
.B1(net137),
.C1(net135),
.Y(net141)
);

sky130_fd_sc_hd__mux4_4 c215(
.A0(net141),
.A1(net14),
.A2(net139),
.A3(net135),
.S0(in27),
.S1(net126),
.X(net142)
);

sky130_fd_sc_hd__nand2b_1 c216(
.A_N(net142),
.B(net674),
.Y(net143)
);

sky130_fd_sc_hd__clkbuf_16 c217(
.A(net627),
.X(net144)
);

sky130_fd_sc_hd__nand3_1 c218(
.A(net11),
.B(net144),
.C(net142),
.Y(net145)
);

sky130_fd_sc_hd__mux4_1 c219(
.A0(net144),
.A1(out35),
.A2(net145),
.A3(net129),
.S0(net139),
.S1(net141),
.X(net146)
);

sky130_fd_sc_hd__or2b_1 c220(
.A(in55),
.B_N(net38),
.X(net147)
);

sky130_fd_sc_hd__nor2_4 c221(
.A(in6),
.B(net43),
.Y(net148)
);

sky130_fd_sc_hd__nand3b_1 c222(
.A_N(net117),
.B(net70),
.C(net42),
.Y(net149)
);

sky130_fd_sc_hd__nand3_2 c223(
.A(net21),
.B(net149),
.C(net127),
.Y(net150)
);

sky130_fd_sc_hd__nor2_4 c224(
.A(net150),
.B(net38),
.Y(net151)
);

sky130_fd_sc_hd__nor3_1 c225(
.A(net30),
.B(net6),
.C(net44),
.Y(net152)
);

sky130_fd_sc_hd__clkinv_8 c226(
.A(net759),
.Y(net153)
);

sky130_fd_sc_hd__and3_2 c227(
.A(net106),
.B(net131),
.C(net38),
.X(net154)
);

sky130_fd_sc_hd__nor2b_4 c228(
.A(net147),
.B_N(net21),
.Y(net155)
);

sky130_fd_sc_hd__nor2b_4 c229(
.A(net36),
.B_N(net154),
.Y(out16)
);

sky130_fd_sc_hd__nor2_2 c230(
.A(net133),
.B(out10),
.Y(net156)
);

sky130_fd_sc_hd__nand3b_4 c231(
.A_N(net156),
.B(net152),
.C(in36),
.Y(net157)
);

sky130_fd_sc_hd__or2b_2 c232(
.A(net44),
.B_N(net131),
.X(out47)
);

sky130_fd_sc_hd__nand2_1 c233(
.A(in0),
.B(net17),
.Y(net158)
);

sky130_fd_sc_hd__nand2_1 c234(
.A(net38),
.B(net152),
.Y(out56)
);

sky130_fd_sc_hd__nor3b_2 c235(
.A(net153),
.B(net140),
.C_N(net28),
.Y(net159)
);

sky130_fd_sc_hd__and3b_1 c236(
.A_N(net28),
.B(out47),
.C(net6),
.X(net160)
);

sky130_fd_sc_hd__o211ai_1 c237(
.A1(net148),
.A2(out56),
.B1(in26),
.C1(net159),
.Y(net161)
);

sky130_fd_sc_hd__nor3_2 c238(
.A(net155),
.B(net158),
.C(net154),
.Y(net162)
);

sky130_fd_sc_hd__or3_1 c239(
.A(net161),
.B(net140),
.C(net162),
.X(net163)
);

sky130_fd_sc_hd__mux4_1 c240(
.A0(net145),
.A1(net160),
.A2(net162),
.A3(net41),
.S0(in45),
.S1(net147),
.X(net164)
);

sky130_fd_sc_hd__mux4_4 c241(
.A0(net6),
.A1(net162),
.A2(net159),
.A3(net147),
.S0(net44),
.S1(net680),
.X(net165)
);

sky130_fd_sc_hd__nor3_2 c242(
.A(net29),
.B(net58),
.C(net681),
.Y(net166)
);

sky130_fd_sc_hd__nor3_1 c243(
.A(net166),
.B(out16),
.C(in20),
.Y(net167)
);

sky130_fd_sc_hd__nand3_4 c244(
.A(net51),
.B(net127),
.C(net60),
.Y(out55)
);

sky130_fd_sc_hd__and3b_4 c245(
.A_N(net160),
.B(net51),
.C(net163),
.X(out60)
);

sky130_fd_sc_hd__o211a_1 c246(
.A1(net118),
.A2(net138),
.B1(out12),
.C1(net163),
.X(out26)
);

sky130_fd_sc_hd__nand3_1 c247(
.A(net127),
.B(out60),
.C(out12),
.Y(net168)
);

sky130_fd_sc_hd__sdfbbn_2 c248(
.D(net142),
.RESET_B(out35),
.SCD(net168),
.SCE(out12),
.SET_B(net62),
.CLK_N(clk),
.Q(net170),
.Q_N(net169)
);

sky130_fd_sc_hd__or3b_2 c249(
.A(net43),
.B(net58),
.C_N(out60),
.X(out44)
);

sky130_fd_sc_hd__o221ai_2 c250(
.A1(in29),
.A2(net43),
.B1(net29),
.B2(net163),
.C1(net169),
.Y(net171)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c251(
.A(net631),
.X(out4)
);

sky130_fd_sc_hd__clkbuf_4 c252(
.A(net630),
.X(net172)
);

sky130_fd_sc_hd__mux4_4 c253(
.A0(net0),
.A1(net169),
.A2(out60),
.A3(net168),
.S0(out4),
.S1(net51),
.X(net173)
);

sky130_fd_sc_hd__o221ai_1 c254(
.A1(net172),
.A2(net138),
.B1(out60),
.B2(net29),
.C1(net683),
.Y(out17)
);

sky130_fd_sc_hd__o221ai_4 c255(
.A1(net170),
.A2(net163),
.B1(out4),
.B2(out60),
.C1(net682),
.Y(net174)
);

sky130_fd_sc_hd__mux4_1 c256(
.A0(net59),
.A1(net167),
.A2(net160),
.A3(out4),
.S0(out17),
.S1(net58),
.X(net175)
);

sky130_fd_sc_hd__o221ai_4 c257(
.A1(net138),
.A2(net170),
.B1(out17),
.B2(net172),
.C1(out35),
.Y(net176)
);

sky130_fd_sc_hd__mux4_4 c258(
.A0(net163),
.A1(net118),
.A2(net43),
.A3(out17),
.S0(out60),
.S1(net682),
.X(net177)
);

sky130_fd_sc_hd__o221a_1 c259(
.A1(net171),
.A2(net172),
.B1(out4),
.B2(net669),
.C1(net684),
.X(net178)
);

sky130_fd_sc_hd__sdfbbp_1 c260(
.D(net60),
.RESET_B(net168),
.SCD(net163),
.SCE(net670),
.SET_B(net681),
.CLK(clk),
.Q(net179)
);

sky130_fd_sc_hd__mux4_1 c261(
.A0(net178),
.A1(out56),
.A2(out57),
.A3(net62),
.S0(net680),
.S1(net684),
.X(net180)
);

sky130_fd_sc_hd__mux4_1 c262(
.A0(net62),
.A1(net174),
.A2(out4),
.A3(net172),
.S0(net682),
.S1(net684),
.X(net181)
);

sky130_fd_sc_hd__mux4_2 c263(
.A0(net179),
.A1(out38),
.A2(out56),
.A3(net118),
.S0(out47),
.S1(out4),
.X(net182)
);

sky130_fd_sc_hd__nand3_4 c264(
.A(net82),
.B(net73),
.C(net64),
.Y(net183)
);

sky130_fd_sc_hd__and2b_1 c265(
.A_N(net67),
.B(net183),
.X(net184)
);

sky130_fd_sc_hd__or3b_1 c266(
.A(net68),
.B(net184),
.C_N(net183),
.X(net185)
);

sky130_fd_sc_hd__nand2b_2 c267(
.A_N(net69),
.B(net183),
.Y(net186)
);

sky130_fd_sc_hd__nor2_4 c268(
.A(in7),
.B(net64),
.Y(net187)
);

sky130_fd_sc_hd__or2_4 c269(
.A(net186),
.B(net183),
.X(net188)
);

sky130_fd_sc_hd__nand2b_4 c270(
.A_N(net65),
.B(in16),
.Y(net189)
);

sky130_fd_sc_hd__nor2_1 c271(
.A(net185),
.B(net73),
.Y(net190)
);

sky130_fd_sc_hd__nand2b_4 c272(
.A_N(net189),
.B(net183),
.Y(net191)
);

sky130_fd_sc_hd__and3b_1 c273(
.A_N(net189),
.B(net191),
.C(net183),
.X(net192)
);

sky130_fd_sc_hd__or2_1 c274(
.A(net77),
.B(net183),
.X(out40)
);

sky130_fd_sc_hd__and2b_1 c275(
.A_N(net184),
.B(net183),
.X(net193)
);

sky130_fd_sc_hd__or2_1 c276(
.A(net73),
.B(net190),
.X(net194)
);

sky130_fd_sc_hd__nand3_2 c277(
.A(net190),
.B(net186),
.C(net183),
.Y(net195)
);

sky130_fd_sc_hd__nor3_4 c278(
.A(in8),
.B(net75),
.C(net81),
.Y(net196)
);

sky130_fd_sc_hd__o221a_2 c279(
.A1(net186),
.A2(net184),
.B1(net195),
.B2(net185),
.C1(net183),
.X(net197)
);

sky130_fd_sc_hd__nand3b_4 c280(
.A_N(net196),
.B(out40),
.C(net183),
.Y(net198)
);

sky130_fd_sc_hd__nand2_2 c281(
.A(net198),
.B(net192),
.Y(net199)
);

sky130_fd_sc_hd__mux4_2 c282(
.A0(net199),
.A1(net188),
.A2(net196),
.A3(out40),
.S0(net64),
.S1(net77),
.X(net200)
);

sky130_fd_sc_hd__nor3_2 c283(
.A(net187),
.B(net198),
.C(net199),
.Y(net201)
);

sky130_fd_sc_hd__o221ai_1 c284(
.A1(net200),
.A2(net78),
.B1(net201),
.B2(net186),
.C1(net183),
.Y(net202)
);

sky130_fd_sc_hd__mux4_4 c285(
.A0(net201),
.A1(net184),
.A2(net196),
.A3(net200),
.S0(net78),
.S1(net188),
.X(out25)
);

sky130_fd_sc_hd__o211a_1 c286(
.A1(net201),
.A2(net74),
.B1(net77),
.C1(net183),
.X(net203)
);

sky130_fd_sc_hd__nor3b_2 c287(
.A(net102),
.B(net88),
.C_N(net201),
.Y(net204)
);

sky130_fd_sc_hd__nor3_2 c288(
.A(net195),
.B(in24),
.C(net77),
.Y(net205)
);

sky130_fd_sc_hd__or3_1 c289(
.A(net194),
.B(net85),
.C(net188),
.X(net206)
);

sky130_fd_sc_hd__o211a_1 c290(
.A1(net188),
.A2(net96),
.B1(in5),
.C1(net94),
.X(net207)
);

sky130_fd_sc_hd__nor2b_2 c291(
.A(net101),
.B_N(net205),
.Y(net208)
);

sky130_fd_sc_hd__and3_4 c292(
.A(net204),
.B(net207),
.C(net94),
.X(net209)
);

sky130_fd_sc_hd__o211ai_4 c293(
.A1(net205),
.A2(in28),
.B1(net194),
.C1(net207),
.Y(net210)
);

sky130_fd_sc_hd__nor2_1 c294(
.A(net209),
.B(net197),
.Y(net211)
);

sky130_fd_sc_hd__or3_4 c295(
.A(net206),
.B(net84),
.C(net94),
.X(net212)
);

sky130_fd_sc_hd__nor3_1 c296(
.A(net212),
.B(net183),
.C(net207),
.Y(net213)
);

sky130_fd_sc_hd__o211ai_2 c297(
.A1(net206),
.A2(net191),
.B1(net203),
.C1(net183),
.Y(net214)
);

sky130_fd_sc_hd__o211ai_4 c298(
.A1(net90),
.A2(net203),
.B1(net201),
.C1(net209),
.Y(net215)
);

sky130_fd_sc_hd__o211a_1 c299(
.A1(net214),
.A2(net209),
.B1(net213),
.C1(net65),
.X(net216)
);

sky130_fd_sc_hd__and2_1 c300(
.A(net203),
.B(net209),
.X(net217)
);

sky130_fd_sc_hd__mux4_2 c301(
.A0(net212),
.A1(net210),
.A2(net200),
.A3(net94),
.S0(net192),
.S1(net217),
.X(net218)
);

sky130_fd_sc_hd__o211a_4 c302(
.A1(in31),
.A2(net216),
.B1(net217),
.C1(net218),
.X(net219)
);

sky130_fd_sc_hd__nor2b_1 c303(
.A(net217),
.B_N(net213),
.Y(net220)
);

sky130_fd_sc_hd__o211a_2 c304(
.A1(net220),
.A2(net219),
.B1(net94),
.C1(net217),
.X(net221)
);

sky130_fd_sc_hd__mux4_2 c305(
.A0(net221),
.A1(net206),
.A2(net211),
.A3(net209),
.S0(out40),
.S1(net94),
.X(net222)
);

sky130_fd_sc_hd__mux4_2 c306(
.A0(net218),
.A1(net217),
.A2(net220),
.A3(in34),
.S0(net207),
.S1(out41),
.X(out46)
);

sky130_fd_sc_hd__mux4_4 c307(
.A0(net204),
.A1(net221),
.A2(net218),
.A3(net220),
.S0(out46),
.S1(net217),
.X(net223)
);

sky130_fd_sc_hd__and3_1 c308(
.A(net207),
.B(in48),
.C(net67),
.X(net224)
);

sky130_fd_sc_hd__or3b_4 c309(
.A(in49),
.B(net207),
.C_N(in43),
.X(net225)
);

sky130_fd_sc_hd__or3_2 c310(
.A(net110),
.B(net121),
.C(net197),
.X(net226)
);

sky130_fd_sc_hd__o211a_1 c311(
.A1(net99),
.A2(net214),
.B1(in45),
.C1(net225),
.X(net227)
);

sky130_fd_sc_hd__o221a_4 c312(
.A1(in57),
.A2(net120),
.B1(net110),
.B2(net224),
.C1(net111),
.X(net228)
);

sky130_fd_sc_hd__nor3_1 c313(
.A(in43),
.B(net123),
.C(net192),
.Y(net229)
);

sky130_fd_sc_hd__nor3b_1 c314(
.A(net203),
.B(net66),
.C_N(net192),
.Y(net230)
);

sky130_fd_sc_hd__nand3b_1 c315(
.A_N(in50),
.B(net116),
.C(net208),
.Y(net231)
);

sky130_fd_sc_hd__nand3b_1 c316(
.A_N(net121),
.B(net229),
.C(net227),
.Y(net232)
);

sky130_fd_sc_hd__o211a_2 c317(
.A1(net210),
.A2(net192),
.B1(net227),
.C1(in43),
.X(net233)
);

sky130_fd_sc_hd__sdfbbn_1 c318(
.D(net232),
.RESET_B(net219),
.SCD(net124),
.SCE(net123),
.SET_B(net203),
.CLK_N(clk),
.Q(out13),
.Q_N(net234)
);

sky130_fd_sc_hd__o211a_4 c319(
.A1(in27),
.A2(net231),
.B1(net234),
.C1(net233),
.X(net235)
);

sky130_fd_sc_hd__o221a_4 c320(
.A1(net227),
.A2(net225),
.B1(net233),
.B2(out13),
.C1(net213),
.X(net236)
);

sky130_fd_sc_hd__sdfrbp_1 c321(
.D(net232),
.RESET_B(net227),
.SCD(net197),
.SCE(net234),
.CLK(clk),
.Q(net238),
.Q_N(net237)
);

sky130_fd_sc_hd__o221ai_2 c322(
.A1(in53),
.A2(in39),
.B1(net226),
.B2(out13),
.C1(net225),
.Y(out23)
);

sky130_fd_sc_hd__buf_2 c323(
.A(net763),
.X(net239)
);

sky130_fd_sc_hd__o221ai_1 c324(
.A1(in39),
.A2(out23),
.B1(net227),
.B2(net233),
.C1(net234),
.Y(net240)
);

sky130_fd_sc_hd__mux4_2 c325(
.A0(net231),
.A1(out13),
.A2(out23),
.A3(net235),
.S0(net111),
.S1(out41),
.X(net241)
);

sky130_fd_sc_hd__o221ai_4 c326(
.A1(net96),
.A2(net232),
.B1(in39),
.B2(net239),
.C1(net234),
.Y(net242)
);

sky130_fd_sc_hd__or3b_4 c327(
.A(net240),
.B(out46),
.C_N(net663),
.X(net243)
);

sky130_fd_sc_hd__mux4_4 c328(
.A0(net240),
.A1(net243),
.A2(in61),
.A3(net237),
.S0(out13),
.S1(net663),
.X(net244)
);

sky130_fd_sc_hd__mux4_2 c329(
.A0(net228),
.A1(in20),
.A2(net238),
.A3(net193),
.S0(net243),
.S1(net685),
.X(net245)
);

sky130_fd_sc_hd__and3_4 c330(
.A(in5),
.B(out13),
.C(net126),
.X(net246)
);

sky130_fd_sc_hd__buf_1 c331(
.A(net637),
.X(out22)
);

sky130_fd_sc_hd__sdfrbp_2 c332(
.D(net128),
.RESET_B(net137),
.SCD(net246),
.SCE(in6),
.CLK(clk),
.Q(net248),
.Q_N(net247)
);

sky130_fd_sc_hd__nand2b_1 c333(
.A_N(net229),
.B(net144),
.Y(net249)
);

sky130_fd_sc_hd__clkinv_2 c334(
.A(net636),
.Y(net250)
);

sky130_fd_sc_hd__nor3b_4 c335(
.A(net140),
.B(net248),
.C_N(net19),
.Y(net251)
);

sky130_fd_sc_hd__nand2b_2 c336(
.A_N(net213),
.B(net17),
.Y(net252)
);

sky130_fd_sc_hd__and2_2 c337(
.A(net251),
.B(in43),
.X(net253)
);

sky130_fd_sc_hd__or2_1 c338(
.A(out35),
.B(net674),
.X(net254)
);

sky130_fd_sc_hd__dlygate4sd3_1 c339(
.A(net760),
.X(net255)
);

sky130_fd_sc_hd__mux4_1 c340(
.A0(net255),
.A1(net104),
.A2(net66),
.A3(net216),
.S0(net254),
.S1(out41),
.X(net256)
);

sky130_fd_sc_hd__nor3b_1 c341(
.A(net248),
.B(net253),
.C_N(net254),
.Y(net257)
);

sky130_fd_sc_hd__mux4_4 c342(
.A0(net257),
.A1(out13),
.A2(net236),
.A3(out23),
.S0(net123),
.S1(net126),
.X(net258)
);

sky130_fd_sc_hd__or3_2 c343(
.A(net235),
.B(net111),
.C(net246),
.X(net259)
);

sky130_fd_sc_hd__or3_4 c344(
.A(net236),
.B(net247),
.C(net257),
.X(out33)
);

sky130_fd_sc_hd__o211a_2 c345(
.A1(net254),
.A2(out53),
.B1(out33),
.C1(net252),
.X(net260)
);

sky130_fd_sc_hd__o211a_2 c346(
.A1(net253),
.A2(net260),
.B1(out33),
.C1(net229),
.X(net261)
);

sky130_fd_sc_hd__o211a_2 c347(
.A1(net260),
.A2(net130),
.B1(out33),
.C1(net132),
.X(net262)
);

sky130_fd_sc_hd__o211ai_4 c348(
.A1(net124),
.A2(net253),
.B1(out33),
.C1(net685),
.Y(net263)
);

sky130_fd_sc_hd__mux4_2 c349(
.A0(net246),
.A1(net235),
.A2(net263),
.A3(out10),
.S0(in29),
.S1(out33),
.X(net264)
);

sky130_fd_sc_hd__mux4_1 c350(
.A0(in61),
.A1(net236),
.A2(net263),
.A3(in34),
.S0(out33),
.S1(out24),
.X(net265)
);

sky130_fd_sc_hd__mux4_2 c351(
.A0(net263),
.A1(net213),
.A2(net260),
.A3(out33),
.S0(out24),
.S1(net686),
.X(net266)
);

sky130_fd_sc_hd__or3_1 c352(
.A(net259),
.B(in47),
.C(net158),
.X(net267)
);

sky130_fd_sc_hd__o221ai_1 c353(
.A1(net66),
.A2(out22),
.B1(out23),
.B2(net685),
.C1(out24),
.Y(out2)
);

sky130_fd_sc_hd__nand3_2 c354(
.A(net17),
.B(net149),
.C(net154),
.Y(out14)
);

sky130_fd_sc_hd__and2b_1 c355(
.A_N(net250),
.B(net17),
.X(net268)
);

sky130_fd_sc_hd__o221a_4 c356(
.A1(net31),
.A2(net165),
.B1(out46),
.B2(net162),
.C1(out33),
.X(out30)
);

sky130_fd_sc_hd__nor3b_1 c357(
.A(in2),
.B(net241),
.C_N(in27),
.Y(net269)
);

sky130_fd_sc_hd__buf_4 c358(
.A(out50),
.X(net270)
);

sky130_fd_sc_hd__or3_1 c359(
.A(net42),
.B(net149),
.C(out46),
.X(out48)
);

sky130_fd_sc_hd__nand3b_4 c360(
.A_N(net157),
.B(net154),
.C(net41),
.Y(net271)
);

sky130_fd_sc_hd__nor3_4 c361(
.A(net132),
.B(net140),
.C(in6),
.Y(out9)
);

sky130_fd_sc_hd__nand3_4 c362(
.A(net197),
.B(out24),
.C(net686),
.Y(net272)
);

sky130_fd_sc_hd__clkinv_16 c363(
.A(net666),
.Y(net273)
);

sky130_fd_sc_hd__o211ai_2 c364(
.A1(net273),
.A2(net270),
.B1(net70),
.C1(out2),
.Y(net274)
);

sky130_fd_sc_hd__o221ai_4 c365(
.A1(net26),
.A2(net159),
.B1(net272),
.B2(out28),
.C1(out30),
.Y(net275)
);

sky130_fd_sc_hd__clkbuf_8 c366(
.A(net759),
.X(net276)
);

sky130_fd_sc_hd__or3b_2 c367(
.A(in36),
.B(net270),
.C_N(net276),
.X(net277)
);

sky130_fd_sc_hd__o211a_2 c368(
.A1(net272),
.A2(net277),
.B1(net149),
.C1(net268),
.X(out54)
);

sky130_fd_sc_hd__sdfbbn_2 c369(
.D(net268),
.RESET_B(net277),
.SCD(out54),
.SCE(out30),
.SET_B(out24),
.CLK_N(clk),
.Q(out51),
.Q_N(net278)
);

sky130_fd_sc_hd__mux4_2 c370(
.A0(net277),
.A1(out54),
.A2(net139),
.A3(out51),
.S0(net152),
.S1(net273),
.X(out36)
);

sky130_fd_sc_hd__o211a_2 c371(
.A1(net271),
.A2(net154),
.B1(out54),
.C1(out41),
.X(net279)
);

sky130_fd_sc_hd__mux4_2 c372(
.A0(in47),
.A1(net279),
.A2(out54),
.A3(out47),
.S0(out23),
.S1(net278),
.X(net280)
);

sky130_fd_sc_hd__mux4_1 c373(
.A0(net267),
.A1(net276),
.A2(out13),
.A3(out54),
.S0(net270),
.S1(net688),
.X(net281)
);

sky130_fd_sc_hd__mux4_4 c392(
.A0(net182),
.A1(out60),
.A2(out38),
.A3(out22),
.S0(out5),
.S1(out40),
.X(out49)
);

sky130_fd_sc_hd__mux4_2 c393(
.A0(net50),
.A1(out58),
.A2(out57),
.A3(out33),
.S0(out28),
.S1(out22),
.X(out52)
);

sky130_fd_sc_hd__mux4_2 c394(
.A0(out49),
.A1(out36),
.A2(net50),
.A3(out4),
.S0(net683),
.S1(net684),
.X(net282)
);

sky130_fd_sc_hd__mux4_4 c395(
.A0(out52),
.A1(net50),
.A2(out61),
.X(out59),
.S0(net683),
.S1(out24)
);

sky130_fd_sc_hd__or2_1 c396(
.A(net190),
.B(net77),
.X(net284)
);

sky130_fd_sc_hd__nor3b_4 c397(
.A(net202),
.B(net193),
.C_N(net183),
.Y(net285)
);

sky130_fd_sc_hd__and2b_2 c398(
.A_N(in5),
.B(in2),
.X(net286)
);

sky130_fd_sc_hd__and3_2 c399(
.A(net74),
.B(net199),
.C(net198),
.X(net287)
);

sky130_fd_sc_hd__nand3_1 c400(
.A(net287),
.B(net76),
.C(net285),
.Y(net288)
);

sky130_fd_sc_hd__o211ai_1 c401(
.A1(net286),
.A2(in17),
.B1(net199),
.C1(net288),
.Y(net289)
);

sky130_fd_sc_hd__nor3_1 c402(
.A(net289),
.B(net288),
.C(net191),
.Y(net290)
);

sky130_fd_sc_hd__o211a_1 c403(
.A1(net285),
.A2(net289),
.B1(net288),
.C1(net197),
.X(net291)
);

sky130_fd_sc_hd__or3b_2 c404(
.A(net291),
.B(net290),
.C_N(net286),
.X(net292)
);

sky130_fd_sc_hd__nor3_4 c405(
.A(net285),
.B(net75),
.C(net190),
.Y(net293)
);

sky130_fd_sc_hd__nor2_1 c406(
.A(net288),
.B(net287),
.Y(net294)
);

sky130_fd_sc_hd__nor3_2 c407(
.A(net80),
.B(net78),
.C(net286),
.Y(net295)
);

sky130_fd_sc_hd__o221ai_1 c408(
.A1(net202),
.A2(net293),
.B1(net288),
.B2(net289),
.C1(net294),
.Y(net296)
);

sky130_fd_sc_hd__mux4_1 c409(
.A0(net294),
.A1(net191),
.A2(net296),
.A3(net193),
.S0(net183),
.S1(net287),
.X(net297)
);

sky130_fd_sc_hd__mux4_2 c410(
.A0(net294),
.A1(net291),
.A2(net288),
.A3(net286),
.S0(net287),
.S1(net183),
.X(net298)
);

sky130_fd_sc_hd__mux4_4 c411(
.A0(net298),
.A1(net297),
.A2(net67),
.A3(net286),
.S0(net289),
.S1(net293),
.X(net299)
);

sky130_fd_sc_hd__mux4_1 c412(
.A0(net290),
.A1(net297),
.A2(net298),
.A3(in6),
.S0(net67),
.S1(net293),
.X(net300)
);

sky130_fd_sc_hd__mux4_2 c413(
.A0(net299),
.A1(net300),
.A2(net294),
.A3(net293),
.S0(net288),
.S1(net298),
.X(net301)
);

sky130_fd_sc_hd__mux4_4 c414(
.A0(net287),
.A1(net293),
.A2(net299),
.A3(net292),
.S0(net288),
.S1(net298),
.X(net302)
);

sky130_fd_sc_hd__mux4_4 c415(
.A0(net293),
.A1(net285),
.A2(net298),
.A3(net295),
.S0(net286),
.S1(net691),
.X(net303)
);

sky130_fd_sc_hd__mux4_4 c416(
.A0(net292),
.A1(net298),
.A2(net293),
.A3(net287),
.S0(net286),
.S1(net659),
.X(net304)
);

sky130_fd_sc_hd__mux4_2 c417(
.A0(net300),
.A1(net303),
.A2(net299),
.A3(net298),
.S0(net304),
.S1(net690),
.X(net305)
);

sky130_fd_sc_hd__nor2_4 c418(
.A(net211),
.B(net75),
.Y(net306)
);

sky130_fd_sc_hd__or3b_4 c419(
.A(net77),
.B(net215),
.C_N(in29),
.X(net307)
);

sky130_fd_sc_hd__and2_2 c420(
.A(net307),
.B(net85),
.X(net308)
);

sky130_fd_sc_hd__and2_1 c421(
.A(net75),
.B(net288),
.X(net309)
);

sky130_fd_sc_hd__nor2_2 c422(
.A(net207),
.B(in29),
.Y(net310)
);

sky130_fd_sc_hd__nor3b_2 c423(
.A(net191),
.B(net84),
.C_N(net77),
.Y(net311)
);

sky130_fd_sc_hd__inv_2 c424(
.A(net623),
.Y(net312)
);

sky130_fd_sc_hd__nor2_2 c425(
.A(in10),
.B(net312),
.Y(net313)
);

sky130_fd_sc_hd__clkinv_2 c426(
.A(net623),
.Y(net314)
);

sky130_fd_sc_hd__mux4_1 c427(
.A0(net217),
.A1(net311),
.A2(net215),
.A3(net313),
.S0(net85),
.S1(net691),
.X(net315)
);

sky130_fd_sc_hd__and2_1 c428(
.A(net88),
.B(net208),
.X(net316)
);

sky130_fd_sc_hd__nand2_1 c429(
.A(net310),
.B(net311),
.Y(net317)
);

sky130_fd_sc_hd__and3_2 c430(
.A(net308),
.B(in24),
.C(net312),
.X(net318)
);

sky130_fd_sc_hd__o221a_4 c431(
.A1(in23),
.A2(net314),
.B1(net94),
.B2(net318),
.C1(net304),
.X(net319)
);

sky130_fd_sc_hd__sdfbbp_1 c432(
.D(net312),
.RESET_B(net315),
.SCD(net311),
.SCE(net318),
.SET_B(net671),
.CLK(clk),
.Q(out19),
.Q_N(net320)
);

sky130_fd_sc_hd__o221ai_2 c433(
.A1(net314),
.A2(out19),
.B1(net312),
.B2(net313),
.C1(net316),
.Y(net321)
);

sky130_fd_sc_hd__buf_8 c434(
.A(net761),
.X(net322)
);

sky130_fd_sc_hd__mux4_2 c435(
.A0(net317),
.A1(net312),
.A2(net293),
.A3(in29),
.S0(net316),
.S1(net671),
.X(net323)
);

sky130_fd_sc_hd__mux4_2 c436(
.A0(net318),
.A1(net215),
.A2(net314),
.A3(net311),
.S0(out41),
.X(net324)
);

sky130_fd_sc_hd__o221ai_2 c437(
.A1(in24),
.A2(net321),
.B1(net288),
.B2(net314),
.C1(net671),
.Y(net325)
);

sky130_fd_sc_hd__o221a_4 c438(
.A1(net325),
.A2(net321),
.B1(net215),
.B2(net658),
.C1(net671),
.X(net326)
);

sky130_fd_sc_hd__and3_2 c439(
.A(net325),
.B(net315),
.C(net671),
.X(net327)
);

sky130_fd_sc_hd__o221a_2 c440(
.A1(net326),
.A2(net183),
.B1(in59),
.B2(net234),
.C1(out28),
.X(net328)
);

sky130_fd_sc_hd__o211a_2 c441(
.A1(net214),
.A2(in58),
.B1(net322),
.C1(net671),
.X(net329)
);

sky130_fd_sc_hd__o221ai_2 c442(
.A1(in54),
.A2(net200),
.B1(out25),
.B2(net233),
.C1(in48),
.Y(net330)
);

sky130_fd_sc_hd__o211a_1 c443(
.A1(net330),
.A2(net313),
.B1(net122),
.C1(in48),
.X(net331)
);

sky130_fd_sc_hd__o211ai_4 c444(
.A1(in59),
.A2(net313),
.B1(net297),
.C1(net316),
.Y(net332)
);

sky130_fd_sc_hd__inv_2 c445(
.A(net626),
.Y(net333)
);

sky130_fd_sc_hd__or3b_2 c446(
.A(net331),
.B(net330),
.C_N(net286),
.X(net334)
);

sky130_fd_sc_hd__o221ai_1 c447(
.A1(net329),
.A2(net230),
.B1(net74),
.B2(net334),
.C1(net296),
.Y(net335)
);

sky130_fd_sc_hd__nand3b_4 c448(
.A_N(net230),
.B(net224),
.C(net286),
.Y(out27)
);

sky130_fd_sc_hd__sdfbbn_1 c449(
.D(net225),
.RESET_B(in59),
.SCD(net197),
.SCE(net334),
.SET_B(net671),
.CLK_N(clk),
.Q(net337),
.Q_N(net336)
);

sky130_fd_sc_hd__sdfbbn_2 c450(
.D(net74),
.RESET_B(net337),
.SCD(in59),
.SCE(net318),
.SET_B(net671),
.CLK_N(clk),
.Q(net339),
.Q_N(net338)
);

sky130_fd_sc_hd__mux4_1 c451(
.A0(net238),
.A1(net230),
.A2(in16),
.A3(in59),
.S0(net337),
.S1(net326),
.X(net340)
);

sky130_fd_sc_hd__buf_6 c452(
.A(net625),
.X(net341)
);

sky130_fd_sc_hd__mux4_2 c453(
.A0(net239),
.A1(net341),
.A2(net339),
.A3(net331),
.S0(in48),
.S1(net336),
.X(net342)
);

sky130_fd_sc_hd__mux4_1 c454(
.A0(net332),
.A1(net340),
.A2(net337),
.A3(net315),
.S0(net331),
.S1(net334),
.X(net343)
);

sky130_fd_sc_hd__o221a_1 c455(
.A1(net231),
.A2(net241),
.B1(net200),
.B2(net336),
.C1(net693),
.X(net344)
);

sky130_fd_sc_hd__o221a_2 c456(
.A1(net233),
.A2(net341),
.B1(net333),
.B2(net337),
.C1(net330),
.X(net345)
);

sky130_fd_sc_hd__mux4_2 c457(
.A0(net345),
.A1(net224),
.A2(net336),
.A3(net333),
.S0(net200),
.S1(net693),
.X(net346)
);

sky130_fd_sc_hd__mux4_1 c458(
.A0(net341),
.A1(net346),
.A2(net331),
.A3(net226),
.S0(net336),
.S1(net692),
.X(net347)
);

sky130_fd_sc_hd__mux4_2 c459(
.A0(net340),
.A1(net331),
.A2(net330),
.A3(net332),
.S0(net321),
.S1(net662),
.X(net348)
);

sky130_fd_sc_hd__mux4_4 c460(
.A0(net344),
.A1(net337),
.A2(net315),
.A3(net233),
.S0(net345),
.S1(net694),
.X(net349)
);

sky130_fd_sc_hd__mux4_2 c461(
.A0(net346),
.A1(net344),
.A2(net334),
.A3(out37),
.S0(net694),
.S1(net695),
.X(net350)
);

sky130_fd_sc_hd__and3b_1 c462(
.A_N(net224),
.B(net130),
.C(net694),
.X(net351)
);

sky130_fd_sc_hd__or2b_4 c463(
.A(net122),
.B_N(net686),
.X(out6)
);

sky130_fd_sc_hd__or3b_1 c464(
.A(net208),
.B(net336),
.C_N(net694),
.X(net352)
);

sky130_fd_sc_hd__nor3_2 c465(
.A(net224),
.B(net256),
.C(net687),
.Y(net353)
);

sky130_fd_sc_hd__or2_4 c466(
.A(net252),
.B(net183),
.X(net354)
);

sky130_fd_sc_hd__and2_0 c467(
.A(net130),
.B(in0),
.X(net355)
);

sky130_fd_sc_hd__and2_1 c468(
.A(net337),
.B(net241),
.X(net356)
);

sky130_fd_sc_hd__nor3_1 c469(
.A(net351),
.B(net126),
.C(out28),
.Y(net357)
);

sky130_fd_sc_hd__or3_1 c470(
.A(net256),
.B(net355),
.C(net352),
.X(net358)
);

sky130_fd_sc_hd__o221a_2 c471(
.A1(net358),
.A2(net352),
.B1(net126),
.B2(net354),
.C1(net686),
.X(net359)
);

sky130_fd_sc_hd__buf_2 c472(
.A(net758),
.X(net360)
);

sky130_fd_sc_hd__mux4_1 c473(
.A0(net126),
.A1(net334),
.A2(net19),
.A3(net356),
.S0(net320),
.S1(net657),
.X(net361)
);

sky130_fd_sc_hd__buf_8 c474(
.A(net757),
.X(net362)
);

sky130_fd_sc_hd__inv_6 c475(
.A(net645),
.Y(net363)
);

sky130_fd_sc_hd__and3b_2 c476(
.A_N(net357),
.B(net351),
.C(out10),
.X(net364)
);

sky130_fd_sc_hd__buf_8 c477(
.A(net644),
.X(net365)
);

sky130_fd_sc_hd__inv_8 c478(
.A(net763),
.Y(net366)
);

sky130_fd_sc_hd__nor3_1 c479(
.A(net284),
.B(net362),
.C(net12),
.Y(net367)
);

sky130_fd_sc_hd__mux4_2 c480(
.A0(net359),
.A1(net360),
.A2(net356),
.A3(out6),
.S0(net365),
.S1(net366),
.X(net368)
);

sky130_fd_sc_hd__and3_1 c481(
.A(net258),
.B(net367),
.C(out0),
.X(net369)
);

sky130_fd_sc_hd__mux4_1 c482(
.A0(net365),
.A1(net369),
.A2(net363),
.A3(net358),
.S0(net356),
.S1(net686),
.X(net370)
);

sky130_fd_sc_hd__inv_16 c483(
.A(net761),
.Y(net371)
);

sky130_fd_sc_hd__o221ai_4 c484(
.A1(net293),
.A2(out33),
.B1(net111),
.B2(net154),
.C1(net688),
.Y(net372)
);

sky130_fd_sc_hd__mux4_1 c485(
.A0(net67),
.A1(out35),
.A2(net41),
.A3(out16),
.S0(out27),
.S1(net234),
.X(net373)
);

sky130_fd_sc_hd__mux4_4 c486(
.A0(in48),
.A1(out35),
.A2(net41),
.A3(net658),
.S0(out8),
.S1(net696),
.X(out20)
);

sky130_fd_sc_hd__mux4_2 c487(
.A0(net154),
.A1(net125),
.A2(net315),
.A3(net34),
.S0(out24),
.S1(net689),
.X(net374)
);

sky130_fd_sc_hd__mux4_4 c488(
.A0(net333),
.A1(net125),
.A2(net41),
.A3(net374),
.S0(net315),
.S1(out8),
.X(net375)
);

sky130_fd_sc_hd__mux4_2 c489(
.A0(net279),
.A1(net111),
.A2(out30),
.A3(net315),
.S0(net369),
.S1(in45),
.X(net376)
);

sky130_fd_sc_hd__o221ai_1 c490(
.A1(net372),
.A2(net41),
.B1(out33),
.B2(net34),
.C1(net293),
.Y(net377)
);

sky130_fd_sc_hd__o221a_2 c491(
.A1(net111),
.A2(net41),
.B1(net374),
.B2(net67),
.C1(out20),
.X(net378)
);

sky130_fd_sc_hd__o221a_1 c492(
.A1(net162),
.A2(out9),
.B1(in19),
.B2(net373),
.C1(net673),
.X(net379)
);

sky130_fd_sc_hd__mux4_4 c493(
.A0(out12),
.A1(net34),
.A2(net162),
.A3(net378),
.S0(net673),
.S1(net689),
.X(net380)
);

sky130_fd_sc_hd__mux4_1 c494(
.A0(net315),
.A1(net378),
.A2(out16),
.A3(net279),
.S0(net688),
.S1(net698),
.X(net381)
);

sky130_fd_sc_hd__mux4_2 c495(
.A0(net378),
.A1(net352),
.A2(net334),
.A3(net374),
.S0(net673),
.S1(net688),
.X(net382)
);

sky130_fd_sc_hd__mux4_1 c496(
.A0(net375),
.A1(net159),
.A2(net374),
.A3(net334),
.S0(net378),
.S1(net698),
.X(net383)
);

sky130_fd_sc_hd__mux4_2 c497(
.A0(net162),
.A1(net369),
.A2(out37),
.A3(out30),
.S0(net41),
.S1(net689),
.X(net384)
);

sky130_fd_sc_hd__sdfbbp_1 c498(
.D(net374),
.RESET_B(net378),
.SCD(net346),
.SCE(out32),
.SET_B(net703),
.CLK(clk),
.Q(out21),
.Q_N(net385)
);

sky130_fd_sc_hd__sdfbbn_1 c499(
.D(net373),
.RESET_B(out30),
.SCD(net699),
.SCE(out32),
.SET_B(net703),
.CLK_N(clk),
.Q(out7),
.Q_N(net386)
);

sky130_fd_sc_hd__mux4_4 c500(
.A0(net366),
.A1(net243),
.A2(net374),
.A3(net352),
.S0(out30),
.S1(net703),
.X(net387)
);

sky130_fd_sc_hd__mux4_1 c501(
.A0(in27),
.A1(net386),
.A2(net352),
.A3(net366),
.S0(net700),
.S1(net704),
.X(net388)
);

sky130_fd_sc_hd__sdfbbn_2 c502(
.D(net354),
.RESET_B(net378),
.SCD(net334),
.SCE(net696),
.SET_B(net704),
.CLK_N(clk),
.Q(net390),
.Q_N(net389)
);

sky130_fd_sc_hd__o221a_2 c503(
.A1(net41),
.A2(out22),
.B1(net315),
.B2(net389),
.C1(net702),
.X(out31)
);

sky130_fd_sc_hd__mux4_2 c504(
.A0(net388),
.A1(net390),
.A2(out7),
.A3(net385),
.S0(net688),
.S1(out32),
.X(net391)
);

sky130_fd_sc_hd__mux4_4 c505(
.A0(net352),
.A1(net391),
.A2(out7),
.A3(net389),
.S0(net698),
.S1(net703),
.X(net392)
);

sky130_fd_sc_hd__or2b_1 c528(
.A(net286),
.B_N(net659),
.X(net393)
);

sky130_fd_sc_hd__and2_1 c529(
.A(net298),
.B(net192),
.X(net394)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c530(
.A(net635),
.X(net395)
);

sky130_fd_sc_hd__nand2b_4 c531(
.A_N(net78),
.B(net287),
.Y(net396)
);

sky130_fd_sc_hd__nand3b_4 c532(
.A_N(net393),
.B(net297),
.C(net289),
.Y(net397)
);

sky130_fd_sc_hd__clkinv_16 c533(
.A(net634),
.Y(net398)
);

sky130_fd_sc_hd__and2_1 c534(
.A(net198),
.B(net395),
.X(net399)
);

sky130_fd_sc_hd__inv_6 c535(
.A(net646),
.Y(net400)
);

sky130_fd_sc_hd__nor3b_1 c536(
.A(net400),
.B(net395),
.C_N(net76),
.Y(net401)
);

sky130_fd_sc_hd__nor2_4 c537(
.A(net396),
.B(net286),
.Y(net402)
);

sky130_fd_sc_hd__and2b_2 c538(
.A_N(net399),
.B(net400),
.X(net403)
);

sky130_fd_sc_hd__nor2b_1 c539(
.A(net400),
.B_N(net399),
.Y(net404)
);

sky130_fd_sc_hd__and2b_2 c540(
.A_N(net291),
.B(net404),
.X(net405)
);

sky130_fd_sc_hd__mux4_2 c541(
.A0(net401),
.A1(net405),
.A2(net402),
.A3(net397),
.S0(net193),
.S1(net199),
.X(net406)
);

sky130_fd_sc_hd__nor2b_1 c542(
.A(net398),
.B_N(net661),
.Y(net407)
);

sky130_fd_sc_hd__inv_6 c543(
.A(net646),
.Y(net408)
);

sky130_fd_sc_hd__o211a_2 c544(
.A1(net408),
.A2(net405),
.B1(net401),
.C1(net395),
.X(net409)
);

sky130_fd_sc_hd__clkinv_1 c545(
.A(net648),
.Y(net410)
);

sky130_fd_sc_hd__o221ai_1 c546(
.A1(net289),
.A2(net410),
.B1(net396),
.B2(net395),
.C1(net401),
.Y(net411)
);

sky130_fd_sc_hd__nor2_1 c547(
.A(net407),
.B(net402),
.Y(net412)
);

sky130_fd_sc_hd__o211ai_2 c548(
.A1(net410),
.A2(net399),
.B1(net409),
.C1(net405),
.Y(net413)
);

sky130_fd_sc_hd__sdfrtn_1 c549(
.D(net412),
.RESET_B(net411),
.SCD(net405),
.SCE(net394),
.CLK_N(clk),
.Q(net414)
);

sky130_fd_sc_hd__nand2_1 c550(
.A(net393),
.B(net322),
.Y(net415)
);

sky130_fd_sc_hd__inv_4 c551(
.A(net633),
.Y(net416)
);

sky130_fd_sc_hd__o221a_2 c552(
.A1(net81),
.A2(net416),
.B1(net313),
.B2(net94),
.C1(net296),
.X(net417)
);

sky130_fd_sc_hd__or2_2 c553(
.A(net323),
.B(net81),
.X(net418)
);

sky130_fd_sc_hd__and2_4 c554(
.A(net415),
.B(net418),
.X(net419)
);

sky130_fd_sc_hd__nor3b_2 c555(
.A(net414),
.B(net321),
.C_N(net402),
.Y(net420)
);

sky130_fd_sc_hd__buf_8 c556(
.A(net632),
.X(net421)
);

sky130_fd_sc_hd__o221a_4 c557(
.A1(in17),
.A2(net192),
.B1(net421),
.B2(net219),
.C1(net419),
.X(net422)
);

sky130_fd_sc_hd__o221a_1 c558(
.A1(net402),
.A2(net327),
.B1(net296),
.B2(net94),
.C1(net419),
.X(net423)
);

sky130_fd_sc_hd__and3_1 c559(
.A(net418),
.B(net323),
.C(net419),
.X(net424)
);

sky130_fd_sc_hd__mux4_2 c560(
.A0(net423),
.A1(net417),
.A2(net424),
.A3(out19),
.S0(net402),
.S1(net419),
.X(net425)
);

sky130_fd_sc_hd__clkbuf_8 c561(
.A(net764),
.X(net426)
);

sky130_fd_sc_hd__inv_8 c562(
.A(net647),
.Y(net427)
);

sky130_fd_sc_hd__o221ai_2 c563(
.A1(net420),
.A2(net427),
.B1(net419),
.B2(net316),
.C1(net655),
.Y(net428)
);

sky130_fd_sc_hd__mux4_1 c564(
.A0(net428),
.A1(net75),
.A2(net394),
.A3(net414),
.S0(net415),
.S1(net419),
.X(net429)
);

sky130_fd_sc_hd__o211a_2 c565(
.A1(net306),
.A2(net417),
.B1(net296),
.C1(net419),
.X(net430)
);

sky130_fd_sc_hd__mux4_2 c566(
.A0(net421),
.A1(net420),
.A2(net427),
.A3(net94),
.S0(net422),
.S1(net397),
.X(net431)
);

sky130_fd_sc_hd__mux4_1 c567(
.A0(net422),
.A1(net219),
.A2(net421),
.A3(net419),
.S0(in14),
.S1(net705),
.X(net432)
);

sky130_fd_sc_hd__sdfbbp_1 c568(
.D(net427),
.RESET_B(net423),
.SCD(net424),
.SCE(net419),
.SET_B(net706),
.CLK(clk),
.Q(net434),
.Q_N(net433)
);

sky130_fd_sc_hd__mux4_1 c569(
.A0(net81),
.A1(net306),
.A2(net427),
.A3(net433),
.S0(net419),
.S1(net661),
.X(net435)
);

sky130_fd_sc_hd__sdfbbn_1 c570(
.D(net435),
.RESET_B(net421),
.SCD(net422),
.SCE(net419),
.SET_B(net654),
.CLK_N(clk),
.Q(net437),
.Q_N(net436)
);

sky130_fd_sc_hd__mux4_4 c571(
.A0(net397),
.A1(net435),
.A2(net417),
.A3(net655),
.S0(net705),
.S1(net706),
.X(net438)
);

sky130_fd_sc_hd__inv_2 c572(
.A(net756),
.Y(net439)
);

sky130_fd_sc_hd__buf_12 c573(
.A(net755),
.X(out11)
);

sky130_fd_sc_hd__nor3_1 c574(
.A(net120),
.B(net239),
.C(out11),
.Y(net440)
);

sky130_fd_sc_hd__clkbuf_8 c575(
.A(net762),
.X(net441)
);

sky130_fd_sc_hd__clkinv_16 c576(
.A(net766),
.Y(net442)
);

sky130_fd_sc_hd__o221ai_1 c577(
.A1(in14),
.A2(net419),
.B1(net338),
.B2(net442),
.C1(net120),
.Y(net443)
);

sky130_fd_sc_hd__o221ai_2 c578(
.A1(net219),
.A2(net296),
.B1(net419),
.B2(net66),
.C1(net707),
.Y(net444)
);

sky130_fd_sc_hd__buf_6 c579(
.A(net765),
.X(net445)
);

sky130_fd_sc_hd__sdfbbn_2 c580(
.D(net441),
.RESET_B(net444),
.SCD(net296),
.SCE(net443),
.SET_B(net707),
.CLK_N(clk),
.Q(net447),
.Q_N(net446)
);

sky130_fd_sc_hd__and3b_1 c581(
.A_N(net322),
.B(net216),
.C(net296),
.X(net448)
);

sky130_fd_sc_hd__nor3b_2 c582(
.A(net339),
.B(net445),
.C_N(in58),
.Y(net449)
);

sky130_fd_sc_hd__sdfbbp_1 c583(
.D(net443),
.RESET_B(net339),
.SCD(net445),
.SCE(net320),
.SET_B(net449),
.CLK(clk),
.Q(net451),
.Q_N(net450)
);

sky130_fd_sc_hd__dlygate4sd1_1 c584(
.A(net764),
.X(net452)
);

sky130_fd_sc_hd__nor3_4 c585(
.A(net452),
.B(net322),
.C(net450),
.Y(net453)
);

sky130_fd_sc_hd__nand3b_4 c586(
.A_N(net445),
.B(net240),
.C(net449),
.Y(net454)
);

sky130_fd_sc_hd__mux4_1 c587(
.A0(net321),
.A1(net221),
.A2(net443),
.A3(net120),
.S0(net451),
.S1(out37),
.X(net455)
);

sky130_fd_sc_hd__mux4_1 c588(
.A0(net328),
.A1(net451),
.A2(net449),
.A3(net694),
.S0(net705),
.S1(net707),
.X(net456)
);

sky130_fd_sc_hd__mux4_1 c589(
.A0(net192),
.A1(net451),
.A2(net342),
.A3(net444),
.S0(net403),
.S1(net443),
.X(net457)
);

sky130_fd_sc_hd__o211ai_1 c590(
.A1(net417),
.A2(net453),
.B1(net676),
.C1(net708),
.Y(net458)
);

sky130_fd_sc_hd__o211a_4 c591(
.A1(net453),
.A2(net111),
.B1(net417),
.C1(net449),
.X(net459)
);

sky130_fd_sc_hd__mux4_4 c592(
.A0(out11),
.A1(net444),
.A2(net240),
.A3(net449),
.S0(net709),
.S1(net710),
.X(net460)
);

sky130_fd_sc_hd__sdfbbn_1 c593(
.D(net232),
.RESET_B(net239),
.SCD(net216),
.SCE(net676),
.SET_B(net694),
.CLK_N(clk),
.Q(net462),
.Q_N(net461)
);

sky130_fd_sc_hd__sdfbbn_2 c594(
.D(net369),
.RESET_B(net221),
.SCD(net125),
.SCE(net449),
.SET_B(net694),
.CLK_N(clk),
.Q(net464),
.Q_N(net463)
);

sky130_fd_sc_hd__mux4_2 c595(
.A0(net104),
.A1(out37),
.A2(net111),
.A3(net125),
.S0(net697),
.S1(net707),
.X(net465)
);

sky130_fd_sc_hd__sdfrtp_1 c596(
.D(net448),
.RESET_B(net197),
.SCD(net334),
.SCE(in34),
.CLK(clk),
.Q(net466)
);

sky130_fd_sc_hd__sdfrtp_2 c597(
.D(net286),
.RESET_B(net466),
.SCD(net369),
.SCE(net111),
.CLK(clk),
.Q(net467)
);

sky130_fd_sc_hd__sdfrtp_4 c598(
.D(net459),
.RESET_B(net448),
.SCD(net234),
.SCE(net705),
.CLK(clk),
.Q(net468)
);

sky130_fd_sc_hd__sdfbbp_1 c599(
.D(net356),
.RESET_B(net466),
.SCD(net468),
.SCE(net369),
.SET_B(net707),
.CLK(clk),
.Q(net470),
.Q_N(net469)
);

sky130_fd_sc_hd__sdfbbn_1 c600(
.D(net466),
.RESET_B(net405),
.SCD(net334),
.SCE(net125),
.SET_B(net468),
.CLK_N(clk),
.Q(net472),
.Q_N(net471)
);

sky130_fd_sc_hd__sdfsbp_1 c601(
.D(net468),
.SCD(net357),
.SCE(net440),
.SET_B(net448),
.CLK(clk),
.Q(net474),
.Q_N(net473)
);

sky130_fd_sc_hd__o221a_1 c602(
.A1(net466),
.A2(net469),
.B1(net12),
.B2(net468),
.C1(net705),
.X(net475)
);

sky130_fd_sc_hd__o221a_4 c603(
.A1(net371),
.A2(net358),
.B1(net459),
.B2(net475),
.C1(out0),
.X(net476)
);

sky130_fd_sc_hd__sdfsbp_2 c604(
.D(net474),
.SCD(net475),
.SCE(net243),
.SET_B(in36),
.CLK(clk),
.Q(net478),
.Q_N(net477)
);

sky130_fd_sc_hd__sdfbbn_2 c605(
.D(net475),
.RESET_B(in16),
.SCD(net461),
.SCE(net369),
.SET_B(net458),
.CLK_N(clk),
.Q(out1),
.Q_N(net479)
);

sky130_fd_sc_hd__mux4_2 c606(
.A0(net465),
.A1(net470),
.A2(out37),
.A3(net444),
.S0(net477),
.S1(net320),
.X(net480)
);

sky130_fd_sc_hd__o221ai_4 c607(
.A1(net478),
.A2(net467),
.B1(net473),
.B2(net667),
.C1(net694),
.Y(net481)
);

sky130_fd_sc_hd__mux4_1 c608(
.A0(net363),
.A1(out1),
.A2(in34),
.A3(net241),
.S0(net467),
.S1(net471),
.X(net482)
);

sky130_fd_sc_hd__o221ai_1 c609(
.A1(net362),
.A2(net472),
.B1(net469),
.B2(net468),
.C1(net694),
.Y(net483)
);

sky130_fd_sc_hd__mux4_1 c610(
.A0(net483),
.A1(net405),
.A2(net481),
.A3(net472),
.S0(net705),
.S1(net710),
.X(net484)
);

sky130_fd_sc_hd__o221a_4 c611(
.A1(in58),
.A2(net481),
.B1(net475),
.B2(net234),
.C1(in27),
.X(net485)
);

sky130_fd_sc_hd__o211ai_1 c612(
.A1(net296),
.A2(net485),
.B1(in2),
.C1(net694),
.Y(net486)
);

sky130_fd_sc_hd__mux4_1 c613(
.A0(net470),
.A1(net484),
.A2(net475),
.A3(net668),
.S0(net694),
.S1(net697),
.X(net487)
);

sky130_fd_sc_hd__mux4_2 c614(
.A0(net440),
.A1(net486),
.A2(in36),
.A3(net484),
.S0(net706),
.S1(net712),
.X(net488)
);

sky130_fd_sc_hd__mux4_2 c615(
.A0(net482),
.A1(net484),
.A2(net125),
.A3(net479),
.S0(out0),
.S1(net713),
.X(net489)
);

sky130_fd_sc_hd__mux4_4 c616(
.A0(net379),
.A1(out19),
.A2(net467),
.A3(net295),
.S0(net34),
.S1(net688),
.X(net490)
);

sky130_fd_sc_hd__mux4_1 c617(
.A0(net374),
.A1(net159),
.A2(net34),
.A3(net386),
.S0(in45),
.S1(net703),
.X(net491)
);

sky130_fd_sc_hd__mux4_4 c618(
.A0(net216),
.A1(in29),
.A2(net158),
.A3(out41),
.S0(net688),
.S1(net714),
.X(net492)
);

sky130_fd_sc_hd__mux4_4 c619(
.A0(net12),
.A1(in45),
.A2(out9),
.A3(out19),
.S0(net385),
.S1(out12),
.X(net493)
);

sky130_fd_sc_hd__mux4_1 c620(
.A0(net492),
.A1(out16),
.A2(net493),
.A3(net482),
.S0(net374),
.S1(net706),
.X(net494)
);

sky130_fd_sc_hd__mux4_4 c621(
.A0(net490),
.A1(net158),
.A2(net320),
.A3(net493),
.S0(net688),
.S1(net702),
.X(net495)
);

sky130_fd_sc_hd__mux4_4 c622(
.A0(net495),
.A1(net358),
.A2(net463),
.A3(net491),
.S0(net386),
.S1(net34),
.X(net496)
);

sky130_fd_sc_hd__mux4_1 c623(
.A0(net334),
.A1(net405),
.A2(net358),
.A3(out13),
.S0(net389),
.S1(net715),
.X(net497)
);

sky130_fd_sc_hd__mux4_4 c624(
.A0(net390),
.A1(net34),
.A2(net159),
.A3(net688),
.S0(net706),
.S1(net707),
.X(net498)
);

sky130_fd_sc_hd__mux4_2 c625(
.A0(net243),
.A1(net492),
.A2(out19),
.A3(net390),
.S0(net491),
.S1(net467),
.X(net499)
);

sky130_fd_sc_hd__mux4_2 c626(
.A0(net491),
.A1(net482),
.A2(net479),
.A3(net707),
.S0(net714),
.S1(net715),
.X(net500)
);

sky130_fd_sc_hd__mux4_1 c627(
.A0(net491),
.A1(net482),
.A2(net493),
.A3(net449),
.S0(net159),
.S1(net216),
.X(net501)
);

sky130_fd_sc_hd__mux4_2 c628(
.A0(net464),
.A1(net498),
.A2(net486),
.A3(out16),
.S0(net491),
.S1(net703),
.X(net502)
);

sky130_fd_sc_hd__mux4_2 c629(
.A0(out14),
.A1(net334),
.A2(net385),
.A3(net707),
.S0(net716),
.S1(net718),
.X(net503)
);

sky130_fd_sc_hd__mux4_2 c630(
.A0(net467),
.A1(net493),
.A2(net320),
.A3(net159),
.S0(out10),
.S1(net717),
.X(net504)
);

sky130_fd_sc_hd__mux4_2 c631(
.A0(net444),
.A1(net159),
.A2(net34),
.A3(net493),
.S0(net717),
.S1(net719),
.X(net505)
);

sky130_fd_sc_hd__mux4_1 c632(
.A0(net221),
.A1(net449),
.A2(net504),
.A3(out21),
.S0(net678),
.S1(net716),
.X(net506)
);

sky130_fd_sc_hd__mux4_4 c633(
.A0(net504),
.A1(net491),
.A2(net243),
.A3(net493),
.S0(net677),
.S1(net721),
.X(net507)
);

sky130_fd_sc_hd__mux4_4 c634(
.A0(net449),
.A1(net295),
.A2(out21),
.A3(net491),
.S0(net706),
.S1(net720),
.X(net508)
);

sky130_fd_sc_hd__mux4_1 c635(
.A0(net493),
.A1(net504),
.A2(net358),
.A3(net706),
.S0(net716),
.S1(net720),
.X(net509)
);

sky130_fd_sc_hd__mux4_1 c636(
.A0(net509),
.A1(out16),
.A2(net504),
.A3(out41),
.S0(net679),
.S1(net688),
.X(net510)
);

sky130_fd_sc_hd__mux4_2 c637(
.A0(net392),
.A1(net491),
.A2(net493),
.A3(net706),
.S0(net719),
.S1(net723),
.X(net511)
);

sky130_fd_sc_hd__clkbuf_1 c660(
.A(net768),
.X(net512)
);

sky130_fd_sc_hd__and2b_4 c661(
.A_N(net404),
.B(net512),
.X(net513)
);

sky130_fd_sc_hd__buf_4 c662(
.A(net675),
.X(net514)
);

sky130_fd_sc_hd__or2b_2 c663(
.A(net407),
.B_N(net199),
.X(net515)
);

sky130_fd_sc_hd__dlygate4sd1_1 c664(
.A(net675),
.X(net516)
);

sky130_fd_sc_hd__or2b_1 c665(
.A(net513),
.B_N(net512),
.X(net517)
);

sky130_fd_sc_hd__nor3b_2 c666(
.A(net399),
.B(net516),
.C_N(net70),
.Y(net518)
);

sky130_fd_sc_hd__or2_4 c667(
.A(net199),
.B(net515),
.X(net519)
);

sky130_fd_sc_hd__nand2b_4 c668(
.A_N(in16),
.B(net512),
.Y(net520)
);

sky130_fd_sc_hd__nand3_1 c669(
.A(net519),
.B(net199),
.C(in16),
.Y(net521)
);

sky130_fd_sc_hd__nor2_1 c670(
.A(net516),
.B(net520),
.Y(net522)
);

sky130_fd_sc_hd__mux4_1 c671(
.A0(net518),
.A1(net522),
.A2(net295),
.A3(net513),
.S0(net512),
.S1(net520),
.X(net523)
);

sky130_fd_sc_hd__o221ai_1 c672(
.A1(net64),
.A2(net409),
.B1(net399),
.B2(in6),
.C1(net513),
.Y(net524)
);

sky130_fd_sc_hd__nand3b_2 c673(
.A_N(net522),
.B(net523),
.C(net660),
.Y(net525)
);

sky130_fd_sc_hd__nand3b_4 c674(
.A_N(net515),
.B(net520),
.C(net660),
.Y(net526)
);

sky130_fd_sc_hd__o221ai_2 c675(
.A1(net515),
.A2(net516),
.B1(net513),
.B2(net512),
.C1(net675),
.Y(net527)
);

sky130_fd_sc_hd__and2b_4 c676(
.A_N(net520),
.B(net521),
.X(net528)
);

sky130_fd_sc_hd__o211a_4 c677(
.A1(net526),
.A2(net528),
.B1(net516),
.C1(net66),
.X(net529)
);

sky130_fd_sc_hd__o211a_2 c678(
.A1(net525),
.A2(net287),
.B1(net522),
.C1(net529),
.X(net530)
);

sky130_fd_sc_hd__inv_2 c679(
.A(net767),
.Y(net531)
);

sky130_fd_sc_hd__o221a_4 c680(
.A1(net527),
.A2(net529),
.B1(net531),
.B2(net530),
.C1(net522),
.X(net532)
);

sky130_fd_sc_hd__o221a_2 c681(
.A1(net521),
.A2(net512),
.B1(net522),
.B2(net513),
.C1(net523),
.X(net533)
);

sky130_fd_sc_hd__nand3_4 c682(
.A(net520),
.B(net434),
.C(net215),
.Y(net534)
);

sky130_fd_sc_hd__o221ai_1 c683(
.A1(net416),
.A2(net426),
.B1(net437),
.B2(net534),
.C1(net533),
.Y(net535)
);

sky130_fd_sc_hd__o211a_1 c684(
.A1(net434),
.A2(in29),
.B1(net316),
.C1(net523),
.X(net536)
);

sky130_fd_sc_hd__o211a_4 c685(
.A1(net437),
.A2(net534),
.B1(net70),
.C1(net516),
.X(net537)
);

sky130_fd_sc_hd__nor3b_2 c686(
.A(net94),
.B(net416),
.C_N(net85),
.Y(net538)
);

sky130_fd_sc_hd__nor3b_4 c687(
.A(net288),
.B(net536),
.C_N(net316),
.Y(net539)
);

sky130_fd_sc_hd__nor3b_2 c688(
.A(net537),
.B(net522),
.C_N(net536),
.Y(net540)
);

sky130_fd_sc_hd__sdfstp_1 c689(
.D(net539),
.SCD(net534),
.SCE(net540),
.SET_B(net538),
.CLK(clk),
.Q(net541)
);

sky130_fd_sc_hd__mux4_4 c690(
.A0(net215),
.A1(net541),
.A2(net419),
.A3(net434),
.S0(net534),
.S1(net532),
.X(net542)
);

sky130_fd_sc_hd__buf_8 c691(
.A(net672),
.X(net543)
);

sky130_fd_sc_hd__o211a_4 c692(
.A1(net522),
.A2(net520),
.B1(net200),
.C1(net542),
.X(net544)
);

sky130_fd_sc_hd__or3_4 c693(
.A(net532),
.B(net414),
.C(net531),
.X(net545)
);

sky130_fd_sc_hd__mux4_1 c694(
.A0(net536),
.A1(net512),
.A2(net535),
.A3(net197),
.S0(net433),
.S1(net419),
.X(net546)
);

sky130_fd_sc_hd__mux4_4 c695(
.A0(net85),
.A1(net538),
.A2(net533),
.A3(net541),
.S0(net316),
.S1(net414),
.X(net547)
);

sky130_fd_sc_hd__sdfbbp_1 c696(
.D(net535),
.RESET_B(net546),
.SCD(net94),
.SCE(net531),
.SET_B(net542),
.CLK(clk),
.Q(net549),
.Q_N(net548)
);

sky130_fd_sc_hd__and3_2 c697(
.A(net517),
.B(net215),
.C(net436),
.X(net550)
);

sky130_fd_sc_hd__o221ai_2 c698(
.A1(net514),
.A2(net416),
.B1(net535),
.B2(net316),
.C1(net419),
.Y(net551)
);

sky130_fd_sc_hd__clkbuf_16 c699(
.A(net672),
.X(net552)
);

sky130_fd_sc_hd__mux4_1 c700(
.A0(net543),
.A1(net548),
.A2(net530),
.A3(net516),
.S0(net94),
.S1(net672),
.X(net553)
);

sky130_fd_sc_hd__mux4_2 c701(
.A0(net530),
.A1(net552),
.A2(net546),
.A3(net550),
.S0(in20),
.S1(net551),
.X(net554)
);

sky130_fd_sc_hd__mux4_1 c702(
.A0(net426),
.A1(net531),
.A2(net433),
.A3(net551),
.S0(net316),
.S1(net725),
.X(net555)
);

sky130_fd_sc_hd__mux4_4 c703(
.A0(net516),
.A1(net316),
.A2(net550),
.A3(net548),
.S0(net540),
.S1(net728),
.X(net556)
);

sky130_fd_sc_hd__o221ai_2 c704(
.A1(net98),
.A2(in20),
.B1(net549),
.B2(net316),
.C1(net543),
.Y(net557)
);

sky130_fd_sc_hd__sdfbbn_1 c705(
.D(net419),
.RESET_B(net551),
.SCD(net403),
.SCE(net450),
.SET_B(net183),
.CLK_N(clk),
.Q(net559),
.Q_N(net558)
);

sky130_fd_sc_hd__o211a_4 c706(
.A1(net553),
.A2(net549),
.B1(net513),
.C1(net711),
.X(net560)
);

sky130_fd_sc_hd__mux4_4 c707(
.A0(net451),
.A1(net534),
.A2(net545),
.A3(net346),
.S0(net216),
.S1(net548),
.X(net561)
);

sky130_fd_sc_hd__o221ai_2 c708(
.A1(net316),
.A2(net513),
.B1(net70),
.B2(net515),
.C1(net730),
.Y(net562)
);

sky130_fd_sc_hd__mux4_2 c709(
.A0(in16),
.A1(out37),
.A2(net553),
.A3(net558),
.S0(net550),
.S1(net523),
.X(net563)
);

sky130_fd_sc_hd__sdfbbn_2 c710(
.D(net560),
.RESET_B(net559),
.SCD(net454),
.SCE(net523),
.SET_B(net419),
.CLK_N(clk),
.Q(net565),
.Q_N(net564)
);

sky130_fd_sc_hd__o211a_2 c711(
.A1(net523),
.A2(net98),
.B1(net559),
.C1(net545),
.X(net566)
);

sky130_fd_sc_hd__mux4_2 c712(
.A0(net443),
.A1(net565),
.A2(net513),
.A3(net653),
.S0(net726),
.S1(net729),
.X(net567)
);

sky130_fd_sc_hd__o211a_2 c713(
.A1(net559),
.A2(in36),
.B1(in58),
.C1(out41),
.X(net568)
);

sky130_fd_sc_hd__mux4_2 c714(
.A0(net533),
.A1(net443),
.A2(net316),
.A3(net454),
.S0(net419),
.S1(out41),
.X(net569)
);

sky130_fd_sc_hd__o221ai_4 c715(
.A1(net442),
.A2(net563),
.B1(net403),
.B2(net533),
.C1(net543),
.Y(net570)
);

sky130_fd_sc_hd__mux4_1 c716(
.A0(net557),
.A1(net450),
.A2(net419),
.A3(net553),
.S0(net727),
.S1(net732),
.X(net571)
);

sky130_fd_sc_hd__o221ai_2 c717(
.A1(net512),
.A2(net419),
.B1(net513),
.B2(net564),
.C1(net732),
.Y(net572)
);

sky130_fd_sc_hd__sdfbbp_1 c718(
.D(net562),
.RESET_B(net216),
.SCD(net571),
.SCE(net513),
.SET_B(net733),
.CLK(clk),
.Q(net573)
);

sky130_fd_sc_hd__sdfstp_2 c719(
.D(net454),
.SCD(net447),
.SCE(net98),
.SET_B(net652),
.CLK(clk),
.Q(net574)
);

sky130_fd_sc_hd__mux4_4 c720(
.A0(net573),
.A1(net572),
.A2(net240),
.A3(net419),
.S0(net730),
.S1(net733),
.X(net575)
);

sky130_fd_sc_hd__o221a_4 c721(
.A1(net559),
.A2(net523),
.B1(out41),
.B2(net726),
.C1(net734),
.X(net576)
);

sky130_fd_sc_hd__mux4_2 c722(
.A0(net576),
.A1(net558),
.A2(net515),
.A3(net419),
.S0(net728),
.S1(net734),
.X(net577)
);

sky130_fd_sc_hd__mux4_4 c723(
.A0(net549),
.A1(net577),
.A2(net558),
.A3(net419),
.S0(net346),
.S1(net734),
.X(net578)
);

sky130_fd_sc_hd__sdfstp_4 c724(
.D(net226),
.SCD(net550),
.SCE(net571),
.SET_B(net735),
.CLK(clk),
.Q(net579)
);

sky130_fd_sc_hd__sdfbbn_1 c725(
.D(net568),
.RESET_B(net574),
.SCD(net98),
.SCE(net579),
.SET_B(net571),
.CLK_N(clk),
.Q(net581),
.Q_N(net580)
);

sky130_fd_sc_hd__mux4_4 c726(
.A0(net297),
.A1(net571),
.A2(net579),
.A3(net541),
.S0(net515),
.S1(in45),
.X(net582)
);

sky130_fd_sc_hd__mux4_2 c727(
.A0(in17),
.A1(net551),
.A2(net197),
.A3(in29),
.S0(net579),
.S1(out41),
.X(net583)
);

sky130_fd_sc_hd__mux4_1 c728(
.A0(net579),
.A1(net297),
.A2(net446),
.A3(in36),
.S0(net665),
.S1(net697),
.X(net584)
);

sky130_fd_sc_hd__sdfbbn_2 c729(
.D(net543),
.RESET_B(net240),
.SCD(net346),
.SCE(net458),
.SET_B(net216),
.CLK_N(clk),
.Q(net586),
.Q_N(net585)
);

sky130_fd_sc_hd__mux4_1 c730(
.A0(net197),
.A1(net515),
.A2(net462),
.A3(net458),
.S0(net545),
.S1(net297),
.X(net587)
);

sky130_fd_sc_hd__mux4_4 c731(
.A0(net447),
.A1(net183),
.A2(net19),
.A3(net66),
.S0(net579),
.S1(net697),
.X(net588)
);

sky130_fd_sc_hd__sdfbbp_1 c732(
.D(net125),
.RESET_B(net346),
.SCD(net541),
.SCE(net710),
.SET_B(net714),
.CLK(clk),
.Q(net589)
);

sky130_fd_sc_hd__o221a_4 c733(
.A1(net565),
.A2(net586),
.B1(net515),
.B2(net580),
.C1(out37),
.X(net590)
);

sky130_fd_sc_hd__mux4_2 c734(
.A0(net200),
.A1(in2),
.A2(net241),
.A3(net66),
.S0(net697),
.S1(net737),
.X(net591)
);

sky130_fd_sc_hd__mux4_1 c735(
.A0(net66),
.A1(net534),
.A2(net564),
.A3(net571),
.S0(net579),
.S1(net590),
.X(net592)
);

sky130_fd_sc_hd__o221ai_1 c736(
.A1(net550),
.A2(net545),
.B1(net591),
.B2(net590),
.C1(net346),
.Y(net593)
);

sky130_fd_sc_hd__sdfbbn_1 c737(
.D(net584),
.RESET_B(net590),
.SCD(net403),
.SCE(net241),
.SET_B(in36),
.CLK_N(clk),
.Q(net594)
);

sky130_fd_sc_hd__mux4_1 c738(
.A0(net403),
.A1(net565),
.A2(net590),
.A3(net591),
.S0(net543),
.S1(out41),
.X(net595)
);

sky130_fd_sc_hd__mux4_1 c739(
.A0(net589),
.A1(net545),
.A2(net590),
.A3(net515),
.S0(net679),
.S1(net739),
.X(net596)
);

sky130_fd_sc_hd__mux4_2 c740(
.A0(net588),
.A1(net590),
.A2(net697),
.A3(net736),
.S0(net739),
.S1(net740),
.X(net597)
);

sky130_fd_sc_hd__mux4_1 c741(
.A0(net19),
.A1(net590),
.A2(net515),
.A3(net597),
.S0(net458),
.S1(net739),
.X(net598)
);

sky130_fd_sc_hd__mux4_2 c742(
.A0(net485),
.A1(net585),
.A2(net590),
.A3(in20),
.S0(net738),
.S1(net739),
.X(net599)
);

sky130_fd_sc_hd__mux4_2 c743(
.A0(net599),
.A1(net591),
.A2(net125),
.A3(net403),
.S0(net597),
.S1(net739),
.X(net600)
);

sky130_fd_sc_hd__mux4_2 c744(
.A0(net579),
.A1(net541),
.A2(net346),
.A3(net597),
.S0(net714),
.S1(net742),
.X(net601)
);

sky130_fd_sc_hd__mux4_2 c745(
.A0(net599),
.A1(in27),
.A2(net550),
.A3(net590),
.S0(net741),
.S1(net742),
.X(net602)
);

sky130_fd_sc_hd__mux4_4 c746(
.A0(net594),
.A1(net484),
.A2(net597),
.A3(net739),
.S0(net742),
.S1(net743),
.X(net603)
);

sky130_fd_sc_hd__mux4_4 c747(
.A0(net597),
.A1(net664),
.A2(net739),
.A3(net742),
.S0(net743),
.S1(net744),
.X(net604)
);

sky130_fd_sc_hd__mux4_2 c748(
.A0(net158),
.A1(net34),
.A2(net701),
.A3(net722),
.S0(net731),
.S1(net739),
.X(net605)
);

sky130_fd_sc_hd__mux4_4 c749(
.A0(net581),
.A1(net605),
.A2(net295),
.A3(net597),
.S0(net484),
.S1(net724),
.X(net606)
);

sky130_fd_sc_hd__mux4_1 c750(
.A0(net241),
.A1(net458),
.A2(net216),
.A3(net547),
.S0(in6),
.S1(net701),
.X(net607)
);

sky130_fd_sc_hd__mux4_2 c751(
.A0(net216),
.A1(net597),
.A2(net346),
.A3(net656),
.S0(net739),
.S1(net745),
.X(net608)
);

sky130_fd_sc_hd__mux4_2 c752(
.A0(net458),
.A1(net547),
.A2(net346),
.A3(net702),
.S0(net739),
.S1(net745),
.X(net609)
);

sky130_fd_sc_hd__mux4_1 c753(
.A0(net125),
.A1(net551),
.A2(net158),
.A3(net604),
.S0(net746),
.S1(net749),
.X(net610)
);

sky130_fd_sc_hd__mux4_2 c754(
.A0(net183),
.A1(in27),
.A2(in20),
.A3(net714),
.S0(net746),
.S1(net750),
.X(net611)
);

sky130_fd_sc_hd__mux4_2 c755(
.A0(net602),
.A1(net484),
.A2(net551),
.A3(net711),
.S0(net724),
.S1(net748),
.X(net612)
);

sky130_fd_sc_hd__mux4_1 c756(
.A0(net604),
.A1(net462),
.A2(net295),
.A3(net486),
.S0(net701),
.S1(net751),
.X(net613)
);

sky130_fd_sc_hd__mux4_1 c757(
.A0(net613),
.A1(net346),
.A2(net611),
.A3(net604),
.S0(net486),
.S1(out41),
.X(net614)
);

sky130_fd_sc_hd__mux4_1 c758(
.A0(net34),
.A1(net125),
.A2(net602),
.A3(net748),
.S0(net750),
.S1(net752),
.X(net615)
);

sky130_fd_sc_hd__mux4_2 c759(
.A0(in45),
.A1(net486),
.A2(net724),
.A3(net731),
.S0(net746),
.S1(net750),
.X(net616)
);

sky130_fd_sc_hd__mux4_4 c760(
.A0(net484),
.A1(net125),
.A2(net711),
.A3(net729),
.S0(net747),
.S1(net749),
.X(net617)
);

sky130_fd_sc_hd__mux4_2 c761(
.A0(net405),
.A1(net70),
.A2(net158),
.A3(net34),
.S0(net749),
.S1(net750),
.X(net618)
);

sky130_fd_sc_hd__mux4_1 c762(
.A0(net547),
.A1(net615),
.A2(net616),
.A3(net745),
.S0(net748),
.S1(net750),
.X(net619)
);

sky130_fd_sc_hd__mux4_2 c763(
.A0(net597),
.A1(in58),
.A2(net749),
.A3(net750),
.S0(net753),
.S1(net754),
.X(net620)
);

sky130_fd_sc_hd__mux4_1 c764(
.A0(net295),
.A1(net618),
.A2(net620),
.A3(net604),
.S0(net597),
.S1(net730),
.X(net621)
);

sky130_fd_sc_hd__o221ai_4 merge765(
.A1(net269),
.A2(out30),
.B1(net31),
.B2(net152),
.C1(out2),
.Y(net622)
);

sky130_fd_sc_hd__clkinv_16 merge766(
.A(net762),
.Y(net623)
);

sky130_fd_sc_hd__mux4_2 merge767(
.A0(net342),
.A1(net219),
.A2(in58),
.A3(net84),
.S0(net328),
.S1(net316),
.X(net624)
);

sky130_fd_sc_hd__sdfbbn_2 merge768(
.D(net297),
.RESET_B(net221),
.SCD(net318),
.SCE(net662),
.SET_B(net663),
.CLK_N(clk),
.Q(net626),
.Q_N(net625)
);

sky130_fd_sc_hd__buf_8 merge769(
.A(net760),
.X(net627)
);

sky130_fd_sc_hd__mux4_1 merge770(
.A0(net355),
.A1(net359),
.A2(net224),
.A3(net360),
.S0(net356),
.S1(net284),
.X(net628)
);

sky130_fd_sc_hd__mux4_4 merge771(
.A0(net542),
.A1(net316),
.A2(net539),
.A3(net540),
.S0(net551),
.S1(net436),
.X(net629)
);

sky130_fd_sc_hd__sdfbbp_1 merge772(
.D(net168),
.RESET_B(net60),
.SCD(out44),
.SCE(net58),
.SET_B(net29),
.CLK(clk),
.Q(net631),
.Q_N(net630)
);

sky130_fd_sc_hd__sedfxbp_1 merge773(
.D(net327),
.DE(net304),
.SCD(net394),
.SCE(net419),
.CLK(clk),
.Q(net633),
.Q_N(net632)
);

sky130_fd_sc_hd__sedfxbp_2 merge774(
.D(net76),
.DE(net394),
.SCD(in6),
.SCE(net397),
.CLK(clk),
.Q(net635),
.Q_N(net634)
);

sky130_fd_sc_hd__sdfbbn_1 merge775(
.D(net143),
.RESET_B(net144),
.SCD(net249),
.SCE(net246),
.SET_B(net235),
.CLK_N(clk),
.Q(net637),
.Q_N(net636)
);

sky130_fd_sc_hd__o211ai_1 merge776(
.A1(net397),
.A2(net512),
.B1(net409),
.C1(net297),
.Y(net638)
);

sky130_fd_sc_hd__mux4_2 merge777(
.A0(net274),
.A1(out46),
.A2(net269),
.A3(net151),
.S0(in47),
.S1(out35),
.X(net639)
);

sky130_fd_sc_hd__mux4_1 merge778(
.A0(net10),
.A1(net128),
.A2(net129),
.A3(net137),
.S0(net143),
.S1(net674),
.X(net640)
);

sky130_fd_sc_hd__mux4_1 merge779(
.A0(net367),
.A1(net369),
.A2(net318),
.A3(net316),
.S0(net671),
.S1(net697),
.X(net641)
);

sky130_fd_sc_hd__mux4_1 merge780(
.A0(net313),
.A1(net328),
.A2(net338),
.A3(net311),
.S0(net304),
.S1(net309),
.X(net642)
);

sky130_fd_sc_hd__mux4_1 merge781(
.A0(net227),
.A1(net228),
.A2(net234),
.A3(net353),
.S0(net365),
.S1(net359),
.X(net643)
);

sky130_fd_sc_hd__sdfbbn_2 merge782(
.D(net356),
.RESET_B(net358),
.SCD(net364),
.SCE(in34),
.SET_B(net657),
.CLK_N(clk),
.Q(net645),
.Q_N(net644)
);

sky130_fd_sc_hd__sedfxtp_1 merge783(
.D(net395),
.DE(net397),
.SCD(net303),
.SCE(net401),
.CLK(clk),
.Q(net646)
);

sky130_fd_sc_hd__sdfbbp_1 merge784(
.D(net304),
.RESET_B(net409),
.SCD(net424),
.SCE(net423),
.SET_B(net419),
.CLK(clk),
.Q(net648),
.Q_N(net647)
);

sky130_fd_sc_hd__mux4_1 merge785(
.A0(net420),
.A1(net422),
.A2(net419),
.A3(net430),
.S0(net450),
.S1(net705),
.X(net649)
);

sky130_fd_sc_hd__mux4_2 merge786(
.A0(net439),
.A1(net403),
.A2(net440),
.A3(net193),
.S0(net316),
.S1(net443),
.X(net650)
);

sky130_fd_sc_hd__mux4_1 merge787(
.A0(net287),
.A1(net397),
.A2(net183),
.A3(net529),
.S0(net409),
.S1(net520),
.X(net651)
);

sky130_fd_sc_hd__dfrbp_1 merge788(
.D(net566),
.RESET_B(net570),
.CLK(clk),
.Q(net653),
.Q_N(net652)
);

sky130_fd_sc_hd__dfrbp_2 merge789(
.D(net425),
.RESET_B(net429),
.CLK(clk),
.Q(net655),
.Q_N(net654)
);

sky130_fd_sc_hd__dfrtn_1 merge790(
.D(net222),
.RESET_B(net223),
.CLK_N(clk),
.Q(out41)
);

sky130_fd_sc_hd__dfrtp_1 merge791(
.D(net621),
.RESET_B(net606),
.CLK(clk),
.Q(net656)
);

sky130_fd_sc_hd__dfrtp_2 merge792(
.D(net261),
.RESET_B(net262),
.CLK(clk),
.Q(net657)
);

sky130_fd_sc_hd__dfrtp_4 merge793(
.D(net361),
.RESET_B(net368),
.CLK(clk),
.Q(out0)
);

sky130_fd_sc_hd__dfsbp_1 merge794(
.D(net301),
.SET_B(net305),
.CLK(clk),
.Q(net659),
.Q_N(net658)
);

sky130_fd_sc_hd__dfsbp_2 merge795(
.D(net406),
.SET_B(net413),
.CLK(clk),
.Q(net661),
.Q_N(net660)
);

sky130_fd_sc_hd__dfstp_1 merge796(
.Q(out59),
.SET_B(net282),
.CLK(clk)
);

sky130_fd_sc_hd__dfstp_2 merge797(
.D(net335),
.SET_B(net347),
.CLK(clk),
.Q(net662)
);

sky130_fd_sc_hd__dfstp_4 merge798(
.D(net245),
.SET_B(net242),
.CLK(clk),
.Q(net663)
);

sky130_fd_sc_hd__dlrbn_1 merge799(
.D(net582),
.RESET_B(net583),
.GATE_N(clk),
.Q(net665),
.Q_N(net664)
);

sky130_fd_sc_hd__dlrbn_2 merge800(
.D(net275),
.RESET_B(net622),
.GATE_N(clk),
.Q(out50),
.Q_N(net666)
);

sky130_fd_sc_hd__dlrbp_1 merge801(
.D(net476),
.RESET_B(net480),
.GATE(clk),
.Q(net668),
.Q_N(net667)
);

sky130_fd_sc_hd__dlrbp_2 merge802(
.D(net176),
.RESET_B(net177),
.GATE(clk),
.Q(net670),
.Q_N(net669)
);

sky130_fd_sc_hd__dlrtn_1 merge803(
.Q(net324),
.RESET_B(net319),
.GATE_N(clk)
);

sky130_fd_sc_hd__dlrtn_2 merge804(
.D(net544),
.RESET_B(net629),
.GATE_N(clk),
.Q(net672)
);

sky130_fd_sc_hd__dlrtn_4 merge805(
.D(net377),
.RESET_B(net376),
.GATE_N(clk),
.Q(net673)
);

sky130_fd_sc_hd__dlrtp_1 merge806(
.D(net134),
.RESET_B(net146),
.GATE(clk),
.Q(net674)
);

sky130_fd_sc_hd__dlrtp_2 merge807(
.D(net524),
.RESET_B(net638),
.GATE(clk),
.Q(net675)
);

sky130_fd_sc_hd__dlrtp_4 merge808(
.D(net460),
.RESET_B(net455),
.GATE(clk),
.Q(net676)
);

sky130_fd_sc_hd__edfxbp_1 merge809(
.D(net494),
.DE(net497),
.CLK(clk),
.Q(net678),
.Q_N(net677)
);

sky130_fd_sc_hd__edfxtp_1 merge810(
.D(net593),
.DE(net501),
.CLK(clk),
.Q(net679)
);

sky130_fd_sc_hd__sdlclkp_1 merge811(
.GATE(net181),
.SCE(net180),
.CLK(clk),
.GCLK(out34)
);

sky130_fd_sc_hd__dfxbp_1 s812(
.D(net164),
.CLK(clk),
.Q(net681),
.Q_N(net680)
);

sky130_fd_sc_hd__dfxbp_2 s813(
.D(net173),
.CLK(clk),
.Q(net683),
.Q_N(net682)
);

sky130_fd_sc_hd__dfxtp_1 s814(
.D(net175),
.CLK(clk),
.Q(net684)
);

sky130_fd_sc_hd__dfxtp_2 s815(
.D(net244),
.CLK(clk),
.Q(net685)
);

sky130_fd_sc_hd__dfxtp_4 s816(
.D(net264),
.CLK(clk),
.Q(out24)
);

sky130_fd_sc_hd__dlclkp_1 s817(
.GATE(net265),
.CLK(clk),
.GCLK(net686)
);

sky130_fd_sc_hd__dlclkp_2 s818(
.GATE(net266),
.CLK(clk),
.GCLK(net687)
);

sky130_fd_sc_hd__dlclkp_4 s819(
.GATE(net280),
.CLK(clk),
.GCLK(net688)
);

sky130_fd_sc_hd__dlxbn_1 s820(
.D(net281),
.GATE_N(clk),
.Q(out8),
.Q_N(net689)
);

sky130_fd_sc_hd__dlxbn_2 s821(
.D(net302),
.GATE_N(clk),
.Q(net691),
.Q_N(net690)
);

sky130_fd_sc_hd__dlxbp_1 s822(
.D(net343),
.GATE(clk),
.Q(net693),
.Q_N(net692)
);

sky130_fd_sc_hd__dlxtn_1 s823(
.D(net348),
.GATE_N(clk),
.Q(net694)
);

sky130_fd_sc_hd__dlxtn_2 s824(
.D(net349),
.GATE_N(clk),
.Q(net695)
);

sky130_fd_sc_hd__dlxtn_4 s825(
.D(net350),
.GATE_N(clk),
.Q(net696)
);

sky130_fd_sc_hd__dlxtp_1 s826(
.D(net370),
.GATE(clk),
.Q(net697)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s827(
.D(net380),
.SLEEP_B(clk),
.Q(net698)
);

sky130_fd_sc_hd__dfxbp_1 s828(
.D(net381),
.CLK(clk),
.Q(net700),
.Q_N(net699)
);

sky130_fd_sc_hd__dfxbp_2 s829(
.D(net382),
.CLK(clk),
.Q(net702),
.Q_N(net701)
);

sky130_fd_sc_hd__dfxtp_1 s830(
.D(net383),
.CLK(clk),
.Q(out32)
);

sky130_fd_sc_hd__dfxtp_2 s831(
.D(net384),
.CLK(clk),
.Q(net703)
);

sky130_fd_sc_hd__dfxtp_4 s832(
.D(net387),
.CLK(clk),
.Q(net704)
);

sky130_fd_sc_hd__dlclkp_1 s833(
.GATE(net431),
.CLK(clk),
.GCLK(net705)
);

sky130_fd_sc_hd__dlclkp_2 s834(
.GATE(net432),
.CLK(clk),
.GCLK(net706)
);

sky130_fd_sc_hd__dlclkp_4 s835(
.GATE(net438),
.CLK(clk),
.GCLK(net707)
);

sky130_fd_sc_hd__dlxbn_1 s836(
.D(net456),
.GATE_N(clk),
.Q(net709),
.Q_N(net708)
);

sky130_fd_sc_hd__dlxbn_2 s837(
.D(net457),
.GATE_N(clk),
.Q(net711),
.Q_N(net710)
);

sky130_fd_sc_hd__dlxbp_1 s838(
.D(net487),
.GATE(clk),
.Q(net712)
);

sky130_fd_sc_hd__dlxtn_1 s839(
.D(net488),
.GATE_N(clk),
.Q(net713)
);

sky130_fd_sc_hd__dlxtn_2 s840(
.D(net489),
.GATE_N(clk),
.Q(net714)
);

sky130_fd_sc_hd__dlxtn_4 s841(
.D(net496),
.GATE_N(clk),
.Q(net715)
);

sky130_fd_sc_hd__dlxtp_1 s842(
.D(net499),
.GATE(clk),
.Q(net716)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s843(
.D(net500),
.SLEEP_B(clk),
.Q(net717)
);

sky130_fd_sc_hd__dfxbp_1 s844(
.D(net502),
.CLK(clk),
.Q(net718)
);

sky130_fd_sc_hd__dfxbp_2 s845(
.D(net503),
.CLK(clk),
.Q(net720),
.Q_N(net719)
);

sky130_fd_sc_hd__dfxtp_1 s846(
.D(net505),
.CLK(clk),
.Q(out18)
);

sky130_fd_sc_hd__dfxtp_2 s847(
.D(net506),
.CLK(clk),
.Q(net721)
);

sky130_fd_sc_hd__dfxtp_4 s848(
.D(net507),
.CLK(clk),
.Q(net722)
);

sky130_fd_sc_hd__dlclkp_1 s849(
.GATE(net508),
.CLK(clk),
.GCLK(out15)
);

sky130_fd_sc_hd__dlclkp_2 s850(
.GATE(net510),
.CLK(clk),
.GCLK(net723)
);

sky130_fd_sc_hd__dlclkp_4 s851(
.GATE(net511),
.CLK(clk),
.GCLK(net724)
);

sky130_fd_sc_hd__dlxbn_1 s852(
.D(net554),
.GATE_N(clk),
.Q(net726),
.Q_N(net725)
);

sky130_fd_sc_hd__dlxbn_2 s853(
.D(net555),
.GATE_N(clk),
.Q(net728),
.Q_N(net727)
);

sky130_fd_sc_hd__dlxbp_1 s854(
.D(net556),
.GATE(clk),
.Q(net730),
.Q_N(net729)
);

sky130_fd_sc_hd__dlxtn_1 s855(
.D(net561),
.GATE_N(clk),
.Q(net731)
);

sky130_fd_sc_hd__dlxtn_2 s856(
.D(net567),
.GATE_N(clk),
.Q(net732)
);

sky130_fd_sc_hd__dlxtn_4 s857(
.D(net569),
.GATE_N(clk),
.Q(net733)
);

sky130_fd_sc_hd__dlxtp_1 s858(
.D(net575),
.GATE(clk),
.Q(net734)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s859(
.D(net578),
.SLEEP_B(clk),
.Q(net735)
);

sky130_fd_sc_hd__dfxbp_1 s860(
.D(net587),
.CLK(clk),
.Q(net737),
.Q_N(net736)
);

sky130_fd_sc_hd__dfxbp_2 s861(
.D(net592),
.CLK(clk),
.Q(net738)
);

sky130_fd_sc_hd__dfxtp_1 s862(
.D(net595),
.CLK(clk),
.Q(net739)
);

sky130_fd_sc_hd__dfxtp_2 s863(
.D(net596),
.CLK(clk),
.Q(net740)
);

sky130_fd_sc_hd__dfxtp_4 s864(
.D(net598),
.CLK(clk),
.Q(net741)
);

sky130_fd_sc_hd__dlclkp_1 s865(
.GATE(net600),
.CLK(clk),
.GCLK(net742)
);

sky130_fd_sc_hd__dlclkp_2 s866(
.GATE(net601),
.CLK(clk),
.GCLK(net743)
);

sky130_fd_sc_hd__dlclkp_4 s867(
.GATE(net603),
.CLK(clk),
.GCLK(net744)
);

sky130_fd_sc_hd__dlxbn_1 s868(
.D(net607),
.GATE_N(clk),
.Q(net746),
.Q_N(net745)
);

sky130_fd_sc_hd__dlxbn_2 s869(
.D(net608),
.GATE_N(clk),
.Q(net747)
);

sky130_fd_sc_hd__dlxbp_1 s870(
.D(net609),
.GATE(clk),
.Q(net749),
.Q_N(net748)
);

sky130_fd_sc_hd__dlxtn_1 s871(
.D(net610),
.GATE_N(clk),
.Q(net750)
);

sky130_fd_sc_hd__dlxtn_2 s872(
.D(net612),
.GATE_N(clk),
.Q(net751)
);

sky130_fd_sc_hd__dlxtn_4 s873(
.D(net614),
.GATE_N(clk),
.Q(net752)
);

sky130_fd_sc_hd__dlxtp_1 s874(
.D(net617),
.GATE(clk),
.Q(net753)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s875(
.D(net619),
.SLEEP_B(clk),
.Q(net754)
);

sky130_fd_sc_hd__dfxbp_1 s876(
.D(net624),
.CLK(clk),
.Q(net756),
.Q_N(net755)
);

sky130_fd_sc_hd__dfxbp_2 s877(
.D(net628),
.CLK(clk),
.Q(net758),
.Q_N(net757)
);

sky130_fd_sc_hd__dfxtp_1 s878(
.D(net639),
.CLK(clk),
.Q(net759)
);

sky130_fd_sc_hd__dfxtp_2 s879(
.D(net640),
.CLK(clk),
.Q(net760)
);

sky130_fd_sc_hd__dfxtp_4 s880(
.D(net641),
.CLK(clk),
.Q(net761)
);

sky130_fd_sc_hd__dlclkp_1 s881(
.GATE(net642),
.CLK(clk),
.GCLK(net762)
);

sky130_fd_sc_hd__dlclkp_2 s882(
.GATE(net643),
.CLK(clk),
.GCLK(net763)
);

sky130_fd_sc_hd__dlclkp_4 s883(
.GATE(net649),
.CLK(clk),
.GCLK(net764)
);

sky130_fd_sc_hd__dlxbn_1 s884(
.D(net650),
.GATE_N(clk),
.Q(net766),
.Q_N(net765)
);

sky130_fd_sc_hd__dlxbn_2 s885(
.D(net651),
.GATE_N(clk),
.Q(net768),
.Q_N(net767)
);


endmodule
