module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net945;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net953;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net948;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net949;
 wire net343;
 wire clknet_0_clk;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net937;
 wire net427;
 wire net942;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net943;
 wire net944;
 wire net946;
 wire net947;
 wire net950;
 wire net951;
 wire net952;
 wire net954;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net758;
 wire clknet_1_0__leaf_net758;
 wire clknet_1_1__leaf_net758;
 wire clknet_0_net431;
 wire clknet_1_0__leaf_net431;
 wire clknet_1_1__leaf_net431;
 wire clknet_0_net674;
 wire clknet_1_0__leaf_net674;
 wire clknet_1_1__leaf_net674;
 wire clknet_0_net465;
 wire clknet_1_0__leaf_net465;
 wire clknet_1_1__leaf_net465;
 wire clknet_0_net582;
 wire clknet_1_0__leaf_net582;
 wire clknet_1_1__leaf_net582;
 wire clknet_0_net611;
 wire clknet_1_0__leaf_net611;
 wire clknet_1_1__leaf_net611;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net470;
 wire clknet_1_0__leaf_net470;
 wire clknet_1_1__leaf_net470;
 wire clknet_0_net720;
 wire clknet_1_0__leaf_net720;
 wire clknet_1_1__leaf_net720;
 wire clknet_0_net492;
 wire clknet_1_0__leaf_net492;
 wire clknet_1_1__leaf_net492;
 wire clknet_0_net472;
 wire clknet_1_0__leaf_net472;
 wire clknet_1_1__leaf_net472;
 wire clknet_0_net471;
 wire clknet_1_0__leaf_net471;
 wire clknet_1_1__leaf_net471;
 wire clknet_0_net824;
 wire clknet_1_0__leaf_net824;
 wire clknet_1_1__leaf_net824;
 wire clknet_0_net832;
 wire clknet_1_0__leaf_net832;
 wire clknet_1_1__leaf_net832;
 wire clknet_0_net461;
 wire clknet_1_0__leaf_net461;
 wire clknet_1_1__leaf_net461;
 wire clknet_0_net702;
 wire clknet_1_0__leaf_net702;
 wire clknet_1_1__leaf_net702;
 wire clknet_0_net757;
 wire clknet_1_0__leaf_net757;
 wire clknet_1_1__leaf_net757;
 wire clknet_0_net232;
 wire clknet_1_0__leaf_net232;
 wire clknet_1_1__leaf_net232;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net339;
 wire clknet_1_0__leaf_net339;
 wire clknet_1_1__leaf_net339;
 wire clknet_0_net336;
 wire clknet_1_0__leaf_net336;
 wire clknet_1_1__leaf_net336;
 wire clknet_0_net345;
 wire clknet_1_0__leaf_net345;
 wire clknet_1_1__leaf_net345;
 wire clknet_0_net341;
 wire clknet_1_0__leaf_net341;
 wire clknet_1_1__leaf_net341;
 wire clknet_0_net228;
 wire clknet_1_0__leaf_net228;
 wire clknet_1_1__leaf_net228;
 wire clknet_0_net230;
 wire clknet_1_0__leaf_net230;
 wire clknet_1_1__leaf_net230;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net739;
 wire clknet_1_0__leaf_net739;
 wire clknet_1_1__leaf_net739;
 wire clknet_0_net574;
 wire clknet_1_0__leaf_net574;
 wire clknet_1_1__leaf_net574;
 wire clknet_0_net741;
 wire clknet_1_0__leaf_net741;
 wire clknet_1_1__leaf_net741;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net849;
 wire clknet_1_0__leaf_net849;
 wire clknet_1_1__leaf_net849;
 wire clknet_0_net721;
 wire clknet_1_0__leaf_net721;
 wire clknet_1_1__leaf_net721;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net740;
 wire clknet_1_0__leaf_net740;
 wire clknet_1_1__leaf_net740;
 wire clknet_0_net703;
 wire clknet_1_0__leaf_net703;
 wire clknet_1_1__leaf_net703;
 wire clknet_0_net689;
 wire clknet_1_0__leaf_net689;
 wire clknet_1_1__leaf_net689;
 wire clknet_0_net859;
 wire clknet_1_0__leaf_net859;
 wire clknet_1_1__leaf_net859;
 wire clknet_0_net688;
 wire clknet_1_0__leaf_net688;
 wire clknet_1_1__leaf_net688;
 wire clknet_0_net687;
 wire clknet_1_0__leaf_net687;
 wire clknet_1_1__leaf_net687;
 wire clknet_0_net868;
 wire clknet_1_0__leaf_net868;
 wire clknet_1_1__leaf_net868;
 wire clknet_0_net827;
 wire clknet_1_0__leaf_net827;
 wire clknet_1_1__leaf_net827;
 wire clknet_0_net170;
 wire clknet_1_0__leaf_net170;
 wire clknet_1_1__leaf_net170;
 wire clknet_0_net673;
 wire clknet_1_0__leaf_net673;
 wire clknet_1_1__leaf_net673;
 wire clknet_0_net434;
 wire clknet_1_0__leaf_net434;
 wire clknet_1_1__leaf_net434;
 wire clknet_0_net445;
 wire clknet_1_0__leaf_net445;
 wire clknet_1_1__leaf_net445;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net843;
 wire clknet_1_0__leaf_net843;
 wire clknet_1_1__leaf_net843;
 wire clknet_0_net487;
 wire clknet_1_0__leaf_net487;
 wire clknet_1_1__leaf_net487;
 wire clknet_0_net457;
 wire clknet_1_0__leaf_net457;
 wire clknet_1_1__leaf_net457;
 wire clknet_0_net454;
 wire clknet_1_0__leaf_net454;
 wire clknet_1_1__leaf_net454;
 wire clknet_0_net453;
 wire clknet_1_0__leaf_net453;
 wire clknet_1_1__leaf_net453;
 wire clknet_0_net438;
 wire clknet_1_0__leaf_net438;
 wire clknet_1_1__leaf_net438;
 wire clknet_0_net440;
 wire clknet_1_0__leaf_net440;
 wire clknet_1_1__leaf_net440;
 wire clknet_0_net545;
 wire clknet_1_0__leaf_net545;
 wire clknet_1_1__leaf_net545;
 wire clknet_0_net547;
 wire clknet_1_0__leaf_net547;
 wire clknet_1_1__leaf_net547;
 wire clknet_0_net427;
 wire clknet_1_0__leaf_net427;
 wire clknet_1_1__leaf_net427;
 wire clknet_0_net429;
 wire clknet_1_0__leaf_net429;
 wire clknet_1_1__leaf_net429;
 wire clknet_0_net586;
 wire clknet_1_0__leaf_net586;
 wire clknet_1_1__leaf_net586;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire net227;
 wire net231;
 wire net238;
 wire net342;
 wire net344;
 wire net426;
 wire net428;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;

 sky130_fd_sc_hd__nor3_1 c100 (.A(net3),
    .B(net10),
    .C(net32),
    .Y(net36));
 sky130_fd_sc_hd__or3b_2 c101 (.A(net32),
    .B(net15),
    .C_N(net869),
    .X(net37));
 sky130_fd_sc_hd__a2111oi_2 c102 (.A1(net31),
    .A2(net37),
    .B1(net32),
    .C1(net12),
    .D1(net805),
    .Y(net38));
 sky130_fd_sc_hd__o2111a_2 c103 (.A1(net28),
    .A2(net38),
    .B1(net37),
    .C1(net36),
    .D1(net20),
    .X(net39));
 sky130_fd_sc_hd__nor4b_1 c104 (.A(net35),
    .B(net787),
    .C(net907),
    .D_N(net913),
    .Y(net40));
 sky130_fd_sc_hd__or4_4 c105 (.A(net7),
    .B(net805),
    .C(net907),
    .D(net35),
    .X(net865));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net37),
    .A1(net31),
    .A2(net811),
    .A3(net39),
    .S0(net907),
    .S1(net35),
    .X(net41));
 sky130_fd_sc_hd__mux4_4 c107 (.A0(net15),
    .A1(net41),
    .A2(net40),
    .A3(net27),
    .S0(net37),
    .S1(net908),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net41),
    .A1(net42),
    .A2(net26),
    .A3(net901),
    .S0(net865),
    .S1(net908),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net901),
    .A1(net43),
    .A2(net41),
    .A3(net908),
    .S0(net28),
    .S1(net33),
    .X(net44));
 sky130_fd_sc_hd__nand3b_4 c110 (.A_N(net24),
    .B(net934),
    .C(net31),
    .Y(net45));
 sky130_fd_sc_hd__o2111a_1 c111 (.A1(net17),
    .A2(net865),
    .B1(net31),
    .C1(net934),
    .D1(net45),
    .X(net46));
 sky130_fd_sc_hd__nor2b_1 c112 (.A(net33),
    .B_N(net44),
    .Y(net47));
 sky130_fd_sc_hd__nor2b_1 c113 (.A(net44),
    .B_N(net45),
    .Y(net48));
 sky130_fd_sc_hd__or2b_1 c114 (.A(net46),
    .B_N(net45),
    .X(net49));
 sky130_fd_sc_hd__nor2_1 c115 (.A(net46),
    .B(net815),
    .Y(net50));
 sky130_fd_sc_hd__nor2b_1 c116 (.A(net773),
    .B_N(net45),
    .Y(net51));
 sky130_fd_sc_hd__nand4b_1 c117 (.A_N(net787),
    .B(net869),
    .C(net865),
    .D(net49),
    .Y(net52));
 sky130_fd_sc_hd__nor2_1 c118 (.A(net49),
    .B(net46),
    .Y(net872));
 sky130_fd_sc_hd__nor2_1 c119 (.A(net51),
    .B(net865),
    .Y(net53));
 sky130_fd_sc_hd__buf_2 c120 (.A(net635),
    .X(net861));
 sky130_fd_sc_hd__and2b_1 c121 (.A_N(net45),
    .B(net861),
    .X(net839));
 sky130_fd_sc_hd__and2_1 c122 (.A(net50),
    .B(net1026),
    .X(net54));
 sky130_fd_sc_hd__nand3b_1 c123 (.A_N(net54),
    .B(net861),
    .C(net45),
    .Y(net55));
 sky130_fd_sc_hd__or2b_1 c124 (.A(net55),
    .B_N(net45),
    .X(net862));
 sky130_fd_sc_hd__mux4_2 c125 (.A0(net762),
    .A1(net55),
    .A2(net839),
    .A3(net44),
    .S0(net861),
    .S1(net54),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net796),
    .A1(net862),
    .A2(net31),
    .A3(net1026),
    .S0(net861),
    .S1(net56),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net53),
    .A1(net862),
    .A2(net33),
    .A3(net55),
    .S0(net1026),
    .S1(net861),
    .X(net58));
 sky130_fd_sc_hd__and3b_1 c128 (.A_N(net55),
    .B(net54),
    .C(net680),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net52),
    .A1(net49),
    .A2(net33),
    .A3(net934),
    .S0(net59),
    .S1(net1008),
    .X(net60));
 sky130_fd_sc_hd__a2111oi_1 c130 (.A1(net52),
    .A2(net839),
    .B1(net16),
    .C1(net664),
    .D1(net681),
    .Y(net828));
 sky130_fd_sc_hd__mux4_2 c131 (.A0(net50),
    .A1(net894),
    .A2(net45),
    .A3(net1028),
    .S0(net664),
    .S1(net681),
    .X(net860));
 sky130_fd_sc_hd__or2b_4 c132 (.A(net793),
    .B_N(net766),
    .X(net61));
 sky130_fd_sc_hd__nor2b_4 c133 (.A(net1031),
    .B_N(net933),
    .Y(net62));
 sky130_fd_sc_hd__and4b_2 c134 (.A_N(net61),
    .B(net818),
    .C(net760),
    .D(net815),
    .X(net63));
 sky130_fd_sc_hd__nor2_4 c135 (.A(net765),
    .B(net933),
    .Y(net64));
 sky130_fd_sc_hd__nand2_4 c136 (.A(net63),
    .B(net64),
    .Y(net65));
 sky130_fd_sc_hd__nand2b_2 c137 (.A_N(net760),
    .B(net63),
    .Y(net66));
 sky130_fd_sc_hd__and2_1 c138 (.A(net773),
    .B(net793),
    .X(net67));
 sky130_fd_sc_hd__nor2b_2 c139 (.A(net62),
    .B_N(net61),
    .Y(net68));
 sky130_fd_sc_hd__or2b_4 c140 (.A(net759),
    .B_N(net765),
    .X(net69));
 sky130_fd_sc_hd__or2b_4 c141 (.A(net65),
    .B_N(net64),
    .X(net70));
 sky130_fd_sc_hd__nand2b_2 c142 (.A_N(net818),
    .B(net67),
    .Y(net71));
 sky130_fd_sc_hd__nor2b_1 c143 (.A(net761),
    .B_N(net815),
    .Y(net72));
 sky130_fd_sc_hd__nand2b_1 c144 (.A_N(net67),
    .B(net68),
    .Y(net73));
 sky130_fd_sc_hd__nand4_4 c145 (.A(net71),
    .B(net69),
    .C(net769),
    .D(net935),
    .Y(net74));
 sky130_fd_sc_hd__and2_2 c146 (.A(net69),
    .B(net68),
    .X(net75));
 sky130_fd_sc_hd__and2_4 c147 (.A(net70),
    .B(net73),
    .X(net76));
 sky130_fd_sc_hd__or3_4 c148 (.A(net766),
    .B(net76),
    .C(net74),
    .X(net77));
 sky130_fd_sc_hd__nor4_1 c149 (.A(net65),
    .B(net74),
    .C(net766),
    .D(net935),
    .Y(net78));
 sky130_fd_sc_hd__and3_4 c150 (.A(net76),
    .B(net928),
    .C(net74),
    .X(net79));
 sky130_fd_sc_hd__nor3_2 c151 (.A(net75),
    .B(net72),
    .C(net73),
    .Y(net80));
 sky130_fd_sc_hd__and2b_2 c152 (.A_N(net76),
    .B(net928),
    .X(net81));
 sky130_fd_sc_hd__and2_4 c153 (.A(net80),
    .B(net81),
    .X(net855));
 sky130_fd_sc_hd__nor2_1 c154 (.A(net73),
    .B(net788),
    .Y(net82));
 sky130_fd_sc_hd__or3b_2 c155 (.A(net797),
    .B(net795),
    .C_N(net791),
    .X(net83));
 sky130_fd_sc_hd__and2b_1 c156 (.A_N(net772),
    .B(net774),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c157 (.A0(net786),
    .A1(net79),
    .A2(net775),
    .A3(net780),
    .S0(net789),
    .S1(net785),
    .X(net85));
 sky130_fd_sc_hd__nand2b_1 c158 (.A_N(net76),
    .B(net65),
    .Y(net86));
 sky130_fd_sc_hd__nand2_2 c159 (.A(net933),
    .B(net80),
    .Y(net87));
 sky130_fd_sc_hd__or2_1 c160 (.A(net785),
    .B(net63),
    .X(net88));
 sky130_fd_sc_hd__and3_2 c161 (.A(net86),
    .B(net87),
    .C(net776),
    .X(net89));
 sky130_fd_sc_hd__or2b_4 c162 (.A(net88),
    .B_N(net89),
    .X(net90));
 sky130_fd_sc_hd__and3_4 c163 (.A(net781),
    .B(net85),
    .C(net769),
    .X(net91));
 sky130_fd_sc_hd__nor3_2 c164 (.A(net795),
    .B(net89),
    .C(net71),
    .Y(net92));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net82),
    .A1(net88),
    .A2(net815),
    .A3(net788),
    .S0(net85),
    .S1(net89),
    .X(net93));
 sky130_fd_sc_hd__and2_1 c166 (.A(net344),
    .B(net90),
    .X(net94));
 sky130_fd_sc_hd__mux4_2 c167 (.A0(net86),
    .A1(net62),
    .A2(net770),
    .A3(net780),
    .S0(net77),
    .S1(net785),
    .X(net95));
 sky130_fd_sc_hd__o2111a_1 c168 (.A1(net91),
    .A2(net93),
    .B1(net776),
    .C1(net95),
    .D1(net92),
    .X(net96));
 sky130_fd_sc_hd__nand4b_4 c169 (.A_N(net96),
    .B(net92),
    .C(net89),
    .D(net87),
    .Y(net97));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net97),
    .A1(net92),
    .A2(net93),
    .A3(net89),
    .S0(net95),
    .S1(net73),
    .X(net98));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net794),
    .A1(net97),
    .A2(net98),
    .A3(net775),
    .S0(net70),
    .S1(net781),
    .X(net99));
 sky130_fd_sc_hd__a2111o_2 c172 (.A1(net84),
    .A2(net89),
    .B1(net95),
    .C1(net99),
    .D1(net77),
    .X(net100));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net66),
    .A1(net98),
    .A2(net99),
    .A3(net771),
    .S0(net91),
    .S1(net95),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c174 (.A0(net792),
    .A1(net99),
    .A2(net101),
    .A3(net780),
    .S0(net90),
    .S1(net100),
    .X(net829));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net100),
    .A1(net85),
    .A2(net101),
    .A3(net93),
    .S0(net90),
    .S1(net99),
    .X(net102));
 sky130_fd_sc_hd__or2_1 c176 (.A(net764),
    .B(net83),
    .X(net103));
 sky130_fd_sc_hd__nand3_2 c177 (.A(net802),
    .B(net80),
    .C(net816),
    .Y(net104));
 sky130_fd_sc_hd__and2b_1 c178 (.A_N(net798),
    .B(net1),
    .X(net105));
 sky130_fd_sc_hd__or2_1 c179 (.A(net806),
    .B(net98),
    .X(net106));
 sky130_fd_sc_hd__and2_1 c180 (.A(net789),
    .B(net806),
    .X(net107));
 sky130_fd_sc_hd__a2111oi_4 c181 (.A1(net102),
    .A2(net799),
    .B1(net814),
    .C1(net91),
    .D1(net762),
    .Y(net108));
 sky130_fd_sc_hd__or2b_1 c182 (.A(net67),
    .B_N(net816),
    .X(net109));
 sky130_fd_sc_hd__or2b_4 c183 (.A(net1),
    .B_N(net813),
    .X(net863));
 sky130_fd_sc_hd__or3b_4 c184 (.A(net80),
    .B(net799),
    .C_N(net863),
    .X(net110));
 sky130_fd_sc_hd__a2111oi_1 c185 (.A1(net109),
    .A2(net863),
    .B1(net110),
    .C1(net77),
    .D1(net100),
    .Y(net111));
 sky130_fd_sc_hd__o2111a_4 c186 (.A1(net107),
    .A2(net906),
    .B1(net77),
    .C1(net863),
    .D1(net87),
    .X(net112));
 sky130_fd_sc_hd__and2_4 c187 (.A(net426),
    .B(net106),
    .X(net113));
 sky130_fd_sc_hd__o2111ai_4 c188 (.A1(net107),
    .A2(net806),
    .B1(net110),
    .C1(net426),
    .D1(net906),
    .Y(net114));
 sky130_fd_sc_hd__a2111o_1 c189 (.A1(net110),
    .A2(net955),
    .B1(net1020),
    .C1(net863),
    .D1(net102),
    .X(net115));
 sky130_fd_sc_hd__nor2b_4 c190 (.A(net112),
    .B_N(net108),
    .Y(net116));
 sky130_fd_sc_hd__or2_1 c191 (.A(net89),
    .B(net116),
    .X(net117));
 sky130_fd_sc_hd__nor2b_4 c192 (.A(net116),
    .B_N(net956),
    .Y(net118));
 sky130_fd_sc_hd__a2111o_4 c193 (.A1(net911),
    .A2(net118),
    .B1(net1),
    .C1(net110),
    .D1(net116),
    .X(net119));
 sky130_fd_sc_hd__a2111o_1 c194 (.A1(net105),
    .A2(net119),
    .B1(net798),
    .C1(net957),
    .D1(net110),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net772),
    .A1(net789),
    .A2(net105),
    .A3(net982),
    .S0(net802),
    .S1(net987),
    .X(net121));
 sky130_fd_sc_hd__a2111o_1 c196 (.A1(net121),
    .A2(net0),
    .B1(net983),
    .C1(net98),
    .D1(net988),
    .X(net122));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net805),
    .A1(net982),
    .A2(net121),
    .A3(net103),
    .S0(net987),
    .X(net123));
 sky130_fd_sc_hd__nand2b_1 c198 (.A_N(net779),
    .B(net892),
    .Y(net124));
 sky130_fd_sc_hd__buf_6 c199 (.A(net1006),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 c200 (.A(net633),
    .X(net125));
 sky130_fd_sc_hd__nand2b_1 c201 (.A_N(net18),
    .B(net63),
    .Y(net126));
 sky130_fd_sc_hd__nand4_2 c202 (.A(net81),
    .B(net18),
    .C(net776),
    .D(net925),
    .Y(net127));
 sky130_fd_sc_hd__and3_4 c203 (.A(net127),
    .B(net16),
    .C(net114),
    .X(net128));
 sky130_fd_sc_hd__or4_2 c204 (.A(net63),
    .B(net929),
    .C(net125),
    .D(net926),
    .X(net129));
 sky130_fd_sc_hd__and2_1 c205 (.A(net125),
    .B(net807),
    .X(net130));
 sky130_fd_sc_hd__nand2_4 c206 (.A(net14),
    .B(net104),
    .Y(net845));
 sky130_fd_sc_hd__and3b_1 c207 (.A_N(net5),
    .B(net426),
    .C(net129),
    .X(net131));
 sky130_fd_sc_hd__nand3_4 c208 (.A(net428),
    .B(net94),
    .C(net128),
    .Y(net132));
 sky130_fd_sc_hd__or3_4 c209 (.A(net131),
    .B(net130),
    .C(net926),
    .X(net133));
 sky130_fd_sc_hd__buf_1 c210 (.A(net1006),
    .X(net134));
 sky130_fd_sc_hd__o2111a_1 c211 (.A1(net130),
    .A2(net128),
    .B1(net816),
    .C1(net929),
    .D1(net773),
    .X(net135));
 sky130_fd_sc_hd__mux4_2 c212 (.A0(net11),
    .A1(net776),
    .A2(net134),
    .A3(net129),
    .S0(net132),
    .S1(net845),
    .X(net852));
 sky130_fd_sc_hd__a2111oi_1 c213 (.A1(net126),
    .A2(net82),
    .B1(net829),
    .C1(net132),
    .D1(net845),
    .Y(net136));
 sky130_fd_sc_hd__nand4_4 c214 (.A(net114),
    .B(net1019),
    .C(net813),
    .D(net133),
    .Y(net137));
 sky130_fd_sc_hd__clkbuf_2 c215 (.A(net632),
    .X(net138));
 sky130_fd_sc_hd__a2111o_1 c216 (.A1(net138),
    .A2(net12),
    .B1(net124),
    .C1(net137),
    .D1(net845),
    .X(net139));
 sky130_fd_sc_hd__and4bb_1 c217 (.A_N(net891),
    .B_N(net137),
    .C(net138),
    .D(net653),
    .X(net140));
 sky130_fd_sc_hd__mux4_4 c218 (.A0(net135),
    .A1(net807),
    .A2(net131),
    .A3(net852),
    .S0(net137),
    .S1(net672),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net138),
    .A1(net891),
    .A2(net118),
    .A3(net137),
    .S0(net1006),
    .S1(net1001),
    .X(net142));
 sky130_fd_sc_hd__nor3b_1 c220 (.A(net816),
    .B(net773),
    .C_N(net865),
    .Y(net143));
 sky130_fd_sc_hd__nor3b_2 c221 (.A(net815),
    .B(net17),
    .C_N(net652),
    .Y(net144));
 sky130_fd_sc_hd__nand2_1 c222 (.A(net12),
    .B(net845),
    .Y(net145));
 sky130_fd_sc_hd__nor3_2 c223 (.A(net344),
    .B(net130),
    .C(net128),
    .Y(net146));
 sky130_fd_sc_hd__nand2b_2 c224 (.A_N(net143),
    .B(net146),
    .Y(net147));
 sky130_fd_sc_hd__nor2_2 c225 (.A(net69),
    .B(net144),
    .Y(net148));
 sky130_fd_sc_hd__nor3_1 c226 (.A(net81),
    .B(net148),
    .C(net128),
    .Y(net149));
 sky130_fd_sc_hd__nor3b_1 c227 (.A(net762),
    .B(net148),
    .C_N(net227),
    .Y(net150));
 sky130_fd_sc_hd__or3_1 c228 (.A(net134),
    .B(net133),
    .C(net128),
    .X(net151));
 sky130_fd_sc_hd__o2111a_1 c229 (.A1(net144),
    .A2(net926),
    .B1(net865),
    .C1(net805),
    .D1(net913),
    .X(net152));
 sky130_fd_sc_hd__or2_1 c230 (.A(net130),
    .B(net863),
    .X(net153));
 sky130_fd_sc_hd__nand2_2 c231 (.A(net149),
    .B(net148),
    .Y(net154));
 sky130_fd_sc_hd__and3_2 c232 (.A(net110),
    .B(net17),
    .C(net153),
    .X(net866));
 sky130_fd_sc_hd__nor3b_2 c233 (.A(net84),
    .B(net933),
    .C_N(net154),
    .Y(net155));
 sky130_fd_sc_hd__a2111oi_1 c234 (.A1(net36),
    .A2(net110),
    .B1(net149),
    .C1(net155),
    .D1(net866),
    .Y(net156));
 sky130_fd_sc_hd__o2111a_1 c235 (.A1(net147),
    .A2(net155),
    .B1(net816),
    .C1(net16),
    .D1(net905),
    .X(net157));
 sky130_fd_sc_hd__o2111a_1 c236 (.A1(net26),
    .A2(net144),
    .B1(net866),
    .C1(net145),
    .D1(net990),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net155),
    .A1(net153),
    .A2(net909),
    .A3(net913),
    .S0(net926),
    .S1(net990),
    .X(net159));
 sky130_fd_sc_hd__and3_2 c238 (.A(net153),
    .B(net852),
    .C(net816),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net153),
    .A1(net160),
    .A2(net845),
    .A3(net144),
    .S0(net110),
    .S1(net100),
    .X(net161));
 sky130_fd_sc_hd__inv_2 c240 (.A(net634),
    .Y(net162));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net162),
    .A1(net866),
    .A2(net160),
    .A3(net143),
    .S0(net913),
    .S1(net158),
    .X(net163));
 sky130_fd_sc_hd__and4b_1 c242 (.A_N(net763),
    .B(net872),
    .C(net148),
    .D(net924),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_1 c243 (.A(net620),
    .X(net875));
 sky130_fd_sc_hd__mux4_4 c244 (.A0(net17),
    .A1(net147),
    .A2(net861),
    .A3(net862),
    .S0(net680),
    .S1(net684),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 c245 (.A(net620),
    .X(net165));
 sky130_fd_sc_hd__nor2b_1 c246 (.A(net148),
    .B_N(net848),
    .Y(net166));
 sky130_fd_sc_hd__nand4b_1 c247 (.A_N(net934),
    .B(net829),
    .C(net148),
    .D(net684),
    .Y(net167));
 sky130_fd_sc_hd__nor2_1 c248 (.A(net16),
    .B(clknet_1_0__leaf_net687),
    .Y(net868));
 sky130_fd_sc_hd__or4b_1 c249 (.A(net165),
    .B(net17),
    .C(net865),
    .D_N(net895),
    .X(net168));
 sky130_fd_sc_hd__sdfrbp_1 c250 (.CLK(clknet_4_10_0_clk),
    .D(net168),
    .RESET_B(net929),
    .SCD(clknet_1_0__leaf_net868),
    .SCE(net784),
    .Q(net831),
    .Q_N(net169));
 sky130_fd_sc_hd__nor4_4 c251 (.A(net45),
    .B(clknet_1_0__leaf_net868),
    .C(net1027),
    .D(net807),
    .Y(net170));
 sky130_fd_sc_hd__or2_1 c252 (.A(net16),
    .B(clknet_1_0__leaf_net170),
    .X(net837));
 sky130_fd_sc_hd__sdfrbp_1 c253 (.CLK(clknet_4_10_0_clk),
    .D(net59),
    .RESET_B(net863),
    .SCD(net148),
    .SCE(clknet_1_1__leaf_net170),
    .Q(net864),
    .Q_N(net171));
 sky130_fd_sc_hd__nor4_1 c254 (.A(net56),
    .B(clknet_1_1__leaf_net170),
    .C(net865),
    .D(net681),
    .Y(net172));
 sky130_fd_sc_hd__a2111o_4 c255 (.A1(net31),
    .A2(clknet_1_1__leaf_net170),
    .B1(net860),
    .C1(net17),
    .D1(net169),
    .X(net173));
 sky130_fd_sc_hd__nand4b_2 c256 (.A_N(net167),
    .B(clknet_1_0__leaf_net170),
    .C(clknet_1_1__leaf_net868),
    .D(net680),
    .Y(net867));
 sky130_fd_sc_hd__nor3_1 c257 (.A(clknet_1_0__leaf_net170),
    .B(net16),
    .C(net773),
    .Y(net825));
 sky130_fd_sc_hd__and4_2 c258 (.A(net1027),
    .B(net839),
    .C(net848),
    .D(net669),
    .X(net844));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net166),
    .A1(net48),
    .A2(net844),
    .A3(net45),
    .S0(net160),
    .S1(net684),
    .X(net174));
 sky130_fd_sc_hd__mux4_2 c260 (.A0(net844),
    .A1(net171),
    .A2(net839),
    .A3(net935),
    .S0(net669),
    .S1(clknet_1_0__leaf_net688),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net59),
    .A1(net862),
    .A2(net31),
    .A3(net844),
    .S0(net684),
    .S1(clknet_1_0__leaf_net688),
    .X(net176));
 sky130_fd_sc_hd__sdfrtn_1 c262 (.CLK_N(clknet_4_10_0_clk),
    .D(net1029),
    .RESET_B(net844),
    .SCD(clknet_1_1__leaf_net688),
    .SCE(clknet_1_0__leaf_net689),
    .Q(net874));
 sky130_fd_sc_hd__mux4_4 c263 (.A0(net874),
    .A1(net763),
    .A2(clknet_1_1__leaf_net868),
    .A3(net863),
    .S0(net678),
    .S1(clknet_1_1__leaf_net689),
    .X(net859));
 sky130_fd_sc_hd__and2_2 c264 (.A(net771),
    .B(net74),
    .X(net177));
 sky130_fd_sc_hd__nand2b_2 c265 (.A_N(net78),
    .B(net177),
    .Y(net178));
 sky130_fd_sc_hd__nor2_2 c266 (.A(net782),
    .B(net770),
    .Y(net179));
 sky130_fd_sc_hd__nor2_2 c267 (.A(net177),
    .B(net815),
    .Y(net180));
 sky130_fd_sc_hd__or3_4 c268 (.A(net820),
    .B(net72),
    .C(net177),
    .X(net181));
 sky130_fd_sc_hd__o2111ai_4 c269 (.A1(net181),
    .A2(net180),
    .B1(net178),
    .C1(net68),
    .D1(net64),
    .Y(net182));
 sky130_fd_sc_hd__or2b_1 c270 (.A(net178),
    .B_N(net182),
    .X(net183));
 sky130_fd_sc_hd__or2_2 c271 (.A(net768),
    .B(net181),
    .X(net184));
 sky130_fd_sc_hd__or3_4 c272 (.A(net1031),
    .B(net75),
    .C(net181),
    .X(net185));
 sky130_fd_sc_hd__and3b_2 c273 (.A_N(net184),
    .B(net68),
    .C(net62),
    .X(net186));
 sky130_fd_sc_hd__nand2b_1 c274 (.A_N(net182),
    .B(net71),
    .Y(net187));
 sky130_fd_sc_hd__nor2b_2 c275 (.A(net179),
    .B_N(net186),
    .Y(net188));
 sky130_fd_sc_hd__nor3b_1 c276 (.A(net188),
    .B(net186),
    .C_N(net782),
    .Y(net189));
 sky130_fd_sc_hd__or3_2 c277 (.A(net180),
    .B(net186),
    .C(net935),
    .X(net190));
 sky130_fd_sc_hd__nand3_2 c278 (.A(net72),
    .B(net769),
    .C(net187),
    .Y(net191));
 sky130_fd_sc_hd__nor3_1 c279 (.A(net190),
    .B(net189),
    .C(net191),
    .Y(net192));
 sky130_fd_sc_hd__and3b_1 c280 (.A_N(net192),
    .B(net184),
    .C(net180),
    .X(net193));
 sky130_fd_sc_hd__and3_1 c281 (.A(net187),
    .B(net183),
    .C(net185),
    .X(net194));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net194),
    .A1(net71),
    .A2(net189),
    .A3(net185),
    .S0(net70),
    .S1(net192),
    .X(net195));
 sky130_fd_sc_hd__nor3_1 c283 (.A(net189),
    .B(net188),
    .C(net194),
    .Y(net196));
 sky130_fd_sc_hd__nor3_2 c284 (.A(net782),
    .B(net187),
    .C(net190),
    .Y(net197));
 sky130_fd_sc_hd__nand3b_2 c285 (.A_N(net183),
    .B(net195),
    .C(net197),
    .Y(net198));
 sky130_fd_sc_hd__and2_1 c286 (.A(net99),
    .B(net777),
    .X(net199));
 sky130_fd_sc_hd__and3b_1 c287 (.A_N(net819),
    .B(net185),
    .C(net70),
    .X(net200));
 sky130_fd_sc_hd__or3_2 c288 (.A(net791),
    .B(net70),
    .C(net90),
    .X(net201));
 sky130_fd_sc_hd__or3b_1 c289 (.A(net71),
    .B(net199),
    .C_N(net182),
    .X(net202));
 sky130_fd_sc_hd__nand3b_4 c290 (.A_N(net96),
    .B(net90),
    .C(net933),
    .Y(net203));
 sky130_fd_sc_hd__a2111o_1 c291 (.A1(net197),
    .A2(net184),
    .B1(net90),
    .C1(net776),
    .D1(net933),
    .X(net204));
 sky130_fd_sc_hd__and3_1 c292 (.A(net769),
    .B(net194),
    .C(net99),
    .X(net205));
 sky130_fd_sc_hd__and3_2 c293 (.A(net179),
    .B(net182),
    .C(net87),
    .X(net206));
 sky130_fd_sc_hd__nand3_1 c294 (.A(net70),
    .B(net95),
    .C(net206),
    .Y(net207));
 sky130_fd_sc_hd__or3_4 c295 (.A(net90),
    .B(net202),
    .C(net195),
    .X(net870));
 sky130_fd_sc_hd__a2111oi_4 c296 (.A1(net95),
    .A2(net199),
    .B1(net771),
    .C1(net904),
    .D1(net179),
    .Y(net208));
 sky130_fd_sc_hd__nand3b_1 c297 (.A_N(net204),
    .B(net193),
    .C(net203),
    .Y(net209));
 sky130_fd_sc_hd__or3b_4 c298 (.A(net92),
    .B(net207),
    .C_N(net904),
    .X(net210));
 sky130_fd_sc_hd__or3_1 c299 (.A(net199),
    .B(net208),
    .C(net195),
    .X(net211));
 sky130_fd_sc_hd__or3_2 c300 (.A(net211),
    .B(net205),
    .C(net904),
    .X(net212));
 sky130_fd_sc_hd__and3_1 c301 (.A(net208),
    .B(net204),
    .C(net777),
    .X(net213));
 sky130_fd_sc_hd__mux4_2 c302 (.A0(net178),
    .A1(net213),
    .A2(net209),
    .A3(net92),
    .S0(net206),
    .S1(net904),
    .X(net214));
 sky130_fd_sc_hd__nor3_1 c303 (.A(net202),
    .B(net967),
    .C(net204),
    .Y(net215));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net205),
    .A1(net87),
    .A2(net904),
    .A3(net213),
    .S0(net95),
    .S1(net215),
    .X(net216));
 sky130_fd_sc_hd__mux4_2 c305 (.A0(net215),
    .A1(net194),
    .A2(net212),
    .A3(net179),
    .S0(net214),
    .S1(net211),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net968),
    .A1(net200),
    .A2(net215),
    .A3(net216),
    .S0(net101),
    .S1(net981),
    .X(net218));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net218),
    .A1(net216),
    .A2(net214),
    .A3(net966),
    .S0(net197),
    .S1(net186),
    .X(net219));
 sky130_fd_sc_hd__or4b_4 c308 (.A(net770),
    .B(net113),
    .C(net193),
    .D_N(net91),
    .X(net220));
 sky130_fd_sc_hd__and2b_1 c309 (.A_N(net800),
    .B(net977),
    .X(net221));
 sky130_fd_sc_hd__or2b_1 c310 (.A(net801),
    .B_N(net193),
    .X(net222));
 sky130_fd_sc_hd__or4b_4 c311 (.A(net106),
    .B(net769),
    .C(net206),
    .D_N(net220),
    .X(net223));
 sky130_fd_sc_hd__and4bb_1 c312 (.A_N(net770),
    .B_N(net979),
    .C(net984),
    .D(net115),
    .X(net224));
 sky130_fd_sc_hd__a2111oi_1 c313 (.A1(net769),
    .A2(net788),
    .B1(net91),
    .C1(net984),
    .D1(net979),
    .Y(net225));
 sky130_fd_sc_hd__inv_12 c314 (.A(net663),
    .Y(net821));
 sky130_fd_sc_hd__inv_4 c315 (.A(net662),
    .Y(net226));
 sky130_fd_sc_hd__inv_12 c328_10 (.A(net675),
    .Y(net945));
 sky130_fd_sc_hd__or3b_1 c317 (.A(net200),
    .B(net212),
    .C_N(net944),
    .X(net228));
 sky130_fd_sc_hd__or3b_1 c318 (.A(net980),
    .B(net209),
    .C_N(net226),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net222),
    .A1(net821),
    .A2(net943),
    .A3(net904),
    .S0(net829),
    .S1(net958),
    .X(net230));
 sky130_fd_sc_hd__inv_1 c449_18 (.A(clknet_1_1__leaf_net757),
    .Y(net953));
 sky130_fd_sc_hd__mux4_4 c321 (.A0(net952),
    .A1(net801),
    .A2(net118),
    .A3(net222),
    .S0(net223),
    .S1(net976),
    .X(net232));
 sky130_fd_sc_hd__mux4_2 c322 (.A0(net193),
    .A1(net978),
    .A2(net951),
    .A3(net226),
    .S0(net821),
    .S1(net892),
    .X(net233));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net229),
    .A1(net809),
    .A2(net203),
    .A3(net904),
    .S0(net980),
    .S1(net224),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_16 c324 (.A(net675),
    .X(net235));
 sky130_fd_sc_hd__and3_4 c325 (.A(clknet_1_0__leaf_net232),
    .B(net950),
    .C(net691),
    .X(net849));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(net778),
    .A1(net800),
    .A2(net949),
    .A3(net77),
    .S0(net222),
    .S1(clknet_1_0__leaf_net233),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net235),
    .A1(net959),
    .A2(clknet_1_0__leaf_net230),
    .A3(clknet_1_0__leaf_net849),
    .S0(net805),
    .S1(net691),
    .X(net237));
 sky130_fd_sc_hd__inv_4 c447_13 (.A(net675),
    .Y(net948));
 sky130_fd_sc_hd__mux4_2 c329 (.A0(net87),
    .A1(clknet_1_0__leaf_net232),
    .A2(net118),
    .A3(net206),
    .S0(net62),
    .S1(net663),
    .X(net239));
 sky130_fd_sc_hd__and3b_1 c330 (.A_N(net104),
    .B(net127),
    .C(net820),
    .X(net240));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(net103),
    .A1(net182),
    .A2(net203),
    .A3(net219),
    .S0(net863),
    .S1(net692),
    .X(net241));
 sky130_fd_sc_hd__and3_2 c332 (.A(net813),
    .B(net132),
    .C(net877),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 c333 (.A(net755),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net206),
    .A1(net922),
    .A2(net242),
    .A3(clknet_1_0__leaf_net849),
    .S0(net813),
    .S1(net692),
    .X(net244));
 sky130_fd_sc_hd__o2111a_1 c335 (.A1(net242),
    .A2(net129),
    .B1(net870),
    .C1(net683),
    .D1(net694),
    .X(net245));
 sky130_fd_sc_hd__and3_1 c336 (.A(net799),
    .B(net243),
    .C(net683),
    .X(net246));
 sky130_fd_sc_hd__sdfbbn_1 c337 (.CLK_N(clknet_4_2_0_clk),
    .D(net137),
    .RESET_B(net242),
    .SCD(net845),
    .SCE(net820),
    .SET_B(net694),
    .Q(net248),
    .Q_N(net247));
 sky130_fd_sc_hd__nand3b_1 c338 (.A_N(net118),
    .B(net206),
    .C(net683),
    .Y(net249));
 sky130_fd_sc_hd__or3_2 c339 (.A(net247),
    .B(net693),
    .C(net877),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(net240),
    .A1(net246),
    .A2(net923),
    .A3(net182),
    .S0(net845),
    .S1(net693),
    .X(net251));
 sky130_fd_sc_hd__and3b_1 c341 (.A_N(net251),
    .B(net242),
    .C(net243),
    .X(net252));
 sky130_fd_sc_hd__buf_1 c342 (.A(net755),
    .X(net253));
 sky130_fd_sc_hd__or3_1 c343 (.A(net115),
    .B(net248),
    .C(net246),
    .X(net254));
 sky130_fd_sc_hd__and4_1 c344 (.A(net922),
    .B(net243),
    .C(net246),
    .D(net206),
    .X(net255));
 sky130_fd_sc_hd__a2111o_1 c345 (.A1(net255),
    .A2(net252),
    .B1(net813),
    .C1(net23),
    .D1(net963),
    .X(net256));
 sky130_fd_sc_hd__sdfrtp_4 c346 (.CLK(clknet_4_9_0_clk),
    .D(net245),
    .RESET_B(net905),
    .SCD(clknet_1_0__leaf_net230),
    .SCE(net927),
    .Q(net841));
 sky130_fd_sc_hd__nor4b_4 c347 (.A(net133),
    .B(net841),
    .C(net242),
    .D_N(net1011),
    .Y(net257));
 sky130_fd_sc_hd__and3_1 c348 (.A(net254),
    .B(net775),
    .C(net870),
    .X(net258));
 sky130_fd_sc_hd__or3b_1 c349 (.A(net246),
    .B(net841),
    .C_N(net243),
    .X(net259));
 sky130_fd_sc_hd__nand4_4 c350 (.A(net23),
    .B(net259),
    .C(net922),
    .D(net841),
    .Y(net260));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net94),
    .A1(net248),
    .A2(net820),
    .A3(net260),
    .S0(net137),
    .S1(net995),
    .X(net261));
 sky130_fd_sc_hd__or3b_2 c352 (.A(net250),
    .B(net821),
    .C_N(net841),
    .X(net262));
 sky130_fd_sc_hd__nor3b_2 c353 (.A(net158),
    .B(net100),
    .C_N(net863),
    .Y(net263));
 sky130_fd_sc_hd__nor3b_2 c354 (.A(net146),
    .B(net927),
    .C_N(net26),
    .Y(net264));
 sky130_fd_sc_hd__or3b_2 c355 (.A(net242),
    .B(net262),
    .C_N(net993),
    .X(net265));
 sky130_fd_sc_hd__sdfbbn_1 c356 (.CLK_N(clknet_4_10_0_clk),
    .D(net154),
    .RESET_B(net924),
    .SCD(net934),
    .SCE(clknet_1_1__leaf_net849),
    .SET_B(net929),
    .Q(net873),
    .Q_N(net266));
 sky130_fd_sc_hd__sdfrtp_1 c357 (.CLK(clknet_4_8_0_clk),
    .D(net262),
    .RESET_B(net265),
    .SCD(net250),
    .SCE(net927),
    .Q(net267));
 sky130_fd_sc_hd__and4_1 c358 (.A(net62),
    .B(net905),
    .C(net873),
    .D(net856),
    .X(net268));
 sky130_fd_sc_hd__nor4_1 c359 (.A(net910),
    .B(net262),
    .C(net784),
    .D(net154),
    .Y(net269));
 sky130_fd_sc_hd__sdfbbp_1 c360 (.CLK(clknet_4_10_0_clk),
    .D(net994),
    .RESET_B(net910),
    .SCD(net160),
    .SCE(net262),
    .SET_B(clknet_1_1__leaf_net849),
    .Q(net271),
    .Q_N(net270));
 sky130_fd_sc_hd__sdfrtp_1 c361 (.CLK(clknet_4_9_0_clk),
    .D(net151),
    .RESET_B(net0),
    .SCD(net269),
    .SCE(net263),
    .Q(net272));
 sky130_fd_sc_hd__or3_4 c362 (.A(net271),
    .B(net262),
    .C(net852),
    .X(net273));
 sky130_fd_sc_hd__a2111o_1 c363 (.A1(net934),
    .A2(net150),
    .B1(net152),
    .C1(net268),
    .D1(net273),
    .X(net274));
 sky130_fd_sc_hd__sdfbbn_1 c364 (.CLK_N(clknet_4_8_0_clk),
    .D(net272),
    .RESET_B(net270),
    .SCD(net265),
    .SCE(net219),
    .SET_B(net1009),
    .Q(net276),
    .Q_N(net275));
 sky130_fd_sc_hd__o2111a_1 c365 (.A1(net152),
    .A2(net272),
    .B1(net250),
    .C1(net263),
    .D1(net154),
    .X(net277));
 sky130_fd_sc_hd__sdfbbn_1 c366 (.CLK_N(clknet_4_8_0_clk),
    .D(net226),
    .RESET_B(net160),
    .SCD(net271),
    .SCE(net929),
    .SET_B(net267),
    .Q(net279),
    .Q_N(net278));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net279),
    .A1(net277),
    .A2(net910),
    .A3(net927),
    .S0(net154),
    .S1(net694),
    .X(net280));
 sky130_fd_sc_hd__sdfbbp_1 c368 (.CLK(clknet_4_11_0_clk),
    .D(net276),
    .RESET_B(net271),
    .SCD(net277),
    .SCE(net877),
    .SET_B(net850),
    .Q(net282),
    .Q_N(net281));
 sky130_fd_sc_hd__a2111oi_1 c369 (.A1(net268),
    .A2(net852),
    .B1(net278),
    .C1(net151),
    .D1(net263),
    .Y(net283));
 sky130_fd_sc_hd__sdfbbn_2 c370 (.CLK_N(clknet_4_11_0_clk),
    .D(net277),
    .RESET_B(net886),
    .SCD(net763),
    .SCE(net885),
    .SET_B(net1003),
    .Q(net823),
    .Q_N(net284));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net909),
    .A1(net284),
    .A2(net278),
    .A3(net270),
    .S0(net885),
    .S1(net281),
    .X(net285));
 sky130_fd_sc_hd__mux4_4 c372 (.A0(net275),
    .A1(net279),
    .A2(net284),
    .A3(net885),
    .S1(net685),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net776),
    .A1(net927),
    .A2(net39),
    .A3(net277),
    .S0(net250),
    .S1(net668),
    .X(net287));
 sky130_fd_sc_hd__mux4_4 c392 (.A0(net892),
    .A1(net935),
    .A2(net861),
    .A3(net1027),
    .S0(net147),
    .S1(clknet_1_1__leaf_net868),
    .X(net827));
 sky130_fd_sc_hd__mux4_4 c393 (.A0(net160),
    .A1(net844),
    .A2(clknet_1_0__leaf_net827),
    .A3(net1027),
    .S0(net821),
    .S1(clknet_1_1__leaf_net687),
    .X(net288));
 sky130_fd_sc_hd__mux4_4 c394 (.A0(net807),
    .A1(clknet_1_1__leaf_net827),
    .A2(net865),
    .A3(net860),
    .S0(net871),
    .S1(net850),
    .X(net289));
 sky130_fd_sc_hd__mux4_4 c395 (.A0(net147),
    .A1(clknet_1_0__leaf_net859),
    .A2(clknet_1_0__leaf_net827),
    .A3(net866),
    .S1(net876),
    .X(net290));
 sky130_fd_sc_hd__nor2b_4 c396 (.A(net68),
    .B_N(net75),
    .Y(net291));
 sky130_fd_sc_hd__and3_2 c397 (.A(net768),
    .B(net291),
    .C(net933),
    .X(net292));
 sky130_fd_sc_hd__nor2_2 c398 (.A(net183),
    .B(net292),
    .Y(net293));
 sky130_fd_sc_hd__and2b_1 c399 (.A_N(net293),
    .B(net186),
    .X(net294));
 sky130_fd_sc_hd__nand2b_1 c400 (.A_N(net291),
    .B(net198),
    .Y(net295));
 sky130_fd_sc_hd__nand2_4 c401 (.A(net181),
    .B(net177),
    .Y(net296));
 sky130_fd_sc_hd__nor3b_1 c402 (.A(net192),
    .B(net293),
    .C_N(net186),
    .Y(net297));
 sky130_fd_sc_hd__nor4_1 c403 (.A(net294),
    .B(net183),
    .C(net293),
    .D(net292),
    .Y(net842));
 sky130_fd_sc_hd__nand3b_4 c404 (.A_N(net295),
    .B(net291),
    .C(net918),
    .Y(net298));
 sky130_fd_sc_hd__a2111oi_1 c405 (.A1(net295),
    .A2(net763),
    .B1(net298),
    .C1(net198),
    .D1(net293),
    .Y(net299));
 sky130_fd_sc_hd__or3_1 c406 (.A(net299),
    .B(net66),
    .C(net918),
    .X(net300));
 sky130_fd_sc_hd__or3_4 c407 (.A(net935),
    .B(net768),
    .C(net918),
    .X(net301));
 sky130_fd_sc_hd__nand4b_1 c408 (.A_N(net294),
    .B(net300),
    .C(net291),
    .D(net918),
    .Y(net302));
 sky130_fd_sc_hd__or2b_1 c409 (.A(net302),
    .B_N(net301),
    .X(net303));
 sky130_fd_sc_hd__and3_1 c410 (.A(net917),
    .B(net301),
    .C(net918),
    .X(net304));
 sky130_fd_sc_hd__nand3b_1 c411 (.A_N(net300),
    .B(net917),
    .C(net301),
    .Y(net305));
 sky130_fd_sc_hd__nand3b_4 c412 (.A_N(net293),
    .B(net291),
    .C(net301),
    .Y(net306));
 sky130_fd_sc_hd__nor3b_2 c413 (.A(net198),
    .B(net302),
    .C_N(net306),
    .Y(net307));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net292),
    .A1(net185),
    .A2(net301),
    .A3(net298),
    .S0(net293),
    .S1(net291),
    .X(net308));
 sky130_fd_sc_hd__nand3b_2 c415 (.A_N(net308),
    .B(net768),
    .C(net307),
    .Y(net309));
 sky130_fd_sc_hd__mux4_4 c416 (.A0(net305),
    .A1(net308),
    .A2(net307),
    .A3(net304),
    .S0(net301),
    .S1(net896),
    .X(net310));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net310),
    .A1(net304),
    .A2(net306),
    .A3(net896),
    .S0(net293),
    .S1(net307),
    .X(net311));
 sky130_fd_sc_hd__buf_1 c418 (.A(net677),
    .X(net312));
 sky130_fd_sc_hd__or2_1 c419 (.A(net207),
    .B(net924),
    .X(net313));
 sky130_fd_sc_hd__nor4b_1 c420 (.A(net776),
    .B(net312),
    .C(net774),
    .D_N(net919),
    .Y(net314));
 sky130_fd_sc_hd__or4_4 c421 (.A(net303),
    .B(net201),
    .C(net896),
    .D(net214),
    .X(net315));
 sky130_fd_sc_hd__or3b_1 c422 (.A(net780),
    .B(net315),
    .C_N(net919),
    .X(net316));
 sky130_fd_sc_hd__nand3b_1 c423 (.A_N(net77),
    .B(net904),
    .C(net315),
    .Y(net317));
 sky130_fd_sc_hd__dlygate4sd1_1 c424 (.A(clknet_1_0__leaf_net673),
    .X(net318));
 sky130_fd_sc_hd__sdfbbn_1 c425 (.CLK_N(clknet_4_1_0_clk),
    .D(net924),
    .RESET_B(net219),
    .SCD(net214),
    .SCE(net788),
    .SET_B(net819),
    .Q(net320),
    .Q_N(net319));
 sky130_fd_sc_hd__or3_2 c426 (.A(net214),
    .B(net210),
    .C(net315),
    .X(net321));
 sky130_fd_sc_hd__inv_2 c427 (.A(net677),
    .Y(net322));
 sky130_fd_sc_hd__or3_4 c428 (.A(net180),
    .B(net303),
    .C(net79),
    .X(net323));
 sky130_fd_sc_hd__and3_2 c429 (.A(net305),
    .B(net298),
    .C(net313),
    .X(net324));
 sky130_fd_sc_hd__mux4_2 c430 (.A0(net320),
    .A1(net321),
    .A2(net311),
    .A3(net185),
    .S0(clknet_1_0__leaf_net318),
    .S1(net918),
    .X(net325));
 sky130_fd_sc_hd__or3b_2 c431 (.A(net323),
    .B(net1022),
    .C_N(net319),
    .X(net326));
 sky130_fd_sc_hd__and2_2 c432 (.A(net202),
    .B(net1024),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net186),
    .A1(net296),
    .A2(net203),
    .A3(net323),
    .S0(net321),
    .S1(net918),
    .X(net328));
 sky130_fd_sc_hd__mux4_4 c434 (.A0(net205),
    .A1(net210),
    .A2(net326),
    .A3(net321),
    .S0(net919),
    .S1(net932),
    .X(net329));
 sky130_fd_sc_hd__and4b_1 c435 (.A_N(net326),
    .B(net296),
    .C(net931),
    .D(net698),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net1022),
    .A1(net207),
    .A2(net330),
    .A3(net326),
    .S0(net311),
    .S1(net697),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net321),
    .A1(net330),
    .A2(net212),
    .A3(net1022),
    .S0(net932),
    .S1(net698),
    .X(net332));
 sky130_fd_sc_hd__mux4_4 c438 (.A0(net330),
    .A1(net185),
    .A2(net214),
    .A3(net679),
    .S0(net932),
    .S1(net697),
    .X(net333));
 sky130_fd_sc_hd__mux4_4 c439 (.A0(clknet_1_1__leaf_net318),
    .A1(net326),
    .A2(net320),
    .A3(net330),
    .S1(net679),
    .X(net334));
 sky130_fd_sc_hd__or2_1 c440 (.A(net313),
    .B(net780),
    .X(net335));
 sky130_fd_sc_hd__nor3b_1 c441 (.A(net814),
    .B(net960),
    .C_N(net947),
    .Y(net336));
 sky130_fd_sc_hd__nand2b_1 c442 (.A_N(net312),
    .B(net327),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 c443 (.A(net621),
    .Y(net338));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(net896),
    .A1(clknet_1_0__leaf_net336),
    .A2(clknet_1_1__leaf_net232),
    .A3(net327),
    .S0(net969),
    .S1(net679),
    .X(net339));
 sky130_fd_sc_hd__nand2b_1 c445 (.A_N(net307),
    .B(net323),
    .Y(net340));
 sky130_fd_sc_hd__nor2b_2 c446 (.A(net338),
    .B_N(clknet_1_1__leaf_net336),
    .Y(net341));
 sky130_fd_sc_hd__inv_12 c320_14 (.A(clknet_1_0__leaf_net757),
    .Y(net949));
 sky130_fd_sc_hd__or2b_2 c448 (.A(net335),
    .B_N(net296),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__and2b_4 c450 (.A_N(clknet_1_1__leaf_net336),
    .B(net327),
    .X(net345));
 sky130_fd_sc_hd__nand2b_1 c451 (.A_N(net323),
    .B(net298),
    .Y(net346));
 sky130_fd_sc_hd__sdfbbp_1 c452 (.CLK(clknet_4_1_0_clk),
    .D(net64),
    .RESET_B(net316),
    .SCD(net915),
    .SCE(net690),
    .SET_B(net931),
    .Q(net348),
    .Q_N(net347));
 sky130_fd_sc_hd__inv_4 c453 (.A(net621),
    .Y(net349));
 sky130_fd_sc_hd__or2b_1 c454 (.A(net349),
    .B_N(net971),
    .X(net350));
 sky130_fd_sc_hd__or2_1 c455 (.A(net948),
    .B(net91),
    .X(net351));
 sky130_fd_sc_hd__buf_1 c456 (.A(clknet_1_0__leaf_net758),
    .X(net832));
 sky130_fd_sc_hd__a2111oi_4 c457 (.A1(clknet_1_1__leaf_net233),
    .A2(net323),
    .B1(net338),
    .C1(clknet_1_0__leaf_net341),
    .D1(net690),
    .Y(net352));
 sky130_fd_sc_hd__nand2_1 c458 (.A(net351),
    .B(net954),
    .Y(net353));
 sky130_fd_sc_hd__and2_1 c459 (.A(net340),
    .B(clknet_1_0__leaf_net336),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net354),
    .A1(net224),
    .A2(net915),
    .A3(net0),
    .S0(clknet_1_0__leaf_net832),
    .X(net355));
 sky130_fd_sc_hd__a2111o_2 c461 (.A1(net953),
    .A2(clknet_1_0__leaf_net832),
    .B1(net985),
    .C1(net915),
    .D1(net656),
    .X(net356));
 sky130_fd_sc_hd__and2b_1 c462 (.A_N(net129),
    .B(net915),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 c463 (.A(net630),
    .X(net878));
 sky130_fd_sc_hd__and2_1 c464 (.A(net258),
    .B(net0),
    .X(net358));
 sky130_fd_sc_hd__nand2b_1 c465 (.A_N(net358),
    .B(net91),
    .Y(net359));
 sky130_fd_sc_hd__nand2b_1 c466 (.A_N(net775),
    .B(net23),
    .Y(net834));
 sky130_fd_sc_hd__nor2b_1 c467 (.A(net969),
    .B_N(net670),
    .Y(net360));
 sky130_fd_sc_hd__or3b_2 c468 (.A(net117),
    .B(net127),
    .C_N(net324),
    .X(net361));
 sky130_fd_sc_hd__o2111ai_4 c469 (.A1(net820),
    .A2(net896),
    .B1(net227),
    .C1(net934),
    .D1(net927),
    .Y(net362));
 sky130_fd_sc_hd__and3b_1 c470 (.A_N(net357),
    .B(net132),
    .C(net117),
    .X(net363));
 sky130_fd_sc_hd__mux4_2 c471 (.A0(net363),
    .A1(clknet_1_1__leaf_net232),
    .A2(net962),
    .A3(net311),
    .S0(net889),
    .S1(net927),
    .X(net364));
 sky130_fd_sc_hd__sdfbbn_1 c472 (.CLK_N(clknet_4_3_0_clk),
    .D(net359),
    .RESET_B(net296),
    .SCD(net361),
    .SCE(net845),
    .SET_B(clknet_1_0__leaf_net832),
    .Q(net366),
    .Q_N(net365));
 sky130_fd_sc_hd__inv_12 c473 (.A(net629),
    .Y(net846));
 sky130_fd_sc_hd__nor3_1 c474 (.A(net337),
    .B(net927),
    .C(net258),
    .Y(net367));
 sky130_fd_sc_hd__and3b_1 c475 (.A_N(net346),
    .B(net360),
    .C(net889),
    .X(net830));
 sky130_fd_sc_hd__and3b_1 c476 (.A_N(net182),
    .B(net363),
    .C(clknet_1_0__leaf_net232),
    .X(net368));
 sky130_fd_sc_hd__sdfbbn_1 c477 (.CLK_N(clknet_4_3_0_clk),
    .D(net203),
    .RESET_B(net311),
    .SCD(clknet_1_0__leaf_net230),
    .SCE(net367),
    .SET_B(net929),
    .Q(net370),
    .Q_N(net369));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net961),
    .A1(clknet_1_1__leaf_net339),
    .A2(net23),
    .A3(net986),
    .S0(net878),
    .S1(net203),
    .X(net371));
 sky130_fd_sc_hd__sdfsbp_1 c479 (.CLK(clknet_4_9_0_clk),
    .D(net127),
    .SCD(clknet_1_0__leaf_net368),
    .SCE(net829),
    .SET_B(net889),
    .Q(net373),
    .Q_N(net372));
 sky130_fd_sc_hd__a2111oi_4 c480 (.A1(net370),
    .A2(net846),
    .B1(net358),
    .C1(clknet_1_1__leaf_net232),
    .D1(net889),
    .Y(net374));
 sky130_fd_sc_hd__sdfbbp_1 c481 (.CLK(clknet_4_9_0_clk),
    .D(net132),
    .RESET_B(net182),
    .SCD(clknet_1_0__leaf_net368),
    .SCE(net889),
    .SET_B(net999),
    .Q(net376),
    .Q_N(net375));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net360),
    .A1(net376),
    .A2(net961),
    .A3(net889),
    .S0(net971),
    .S1(clknet_1_0__leaf_net368),
    .X(net377));
 sky130_fd_sc_hd__sdfbbn_1 c483 (.CLK_N(clknet_4_3_0_clk),
    .D(net373),
    .RESET_B(net374),
    .SCD(net375),
    .SCE(net889),
    .SET_B(net369),
    .Q(net379),
    .Q_N(net378));
 sky130_fd_sc_hd__mux4_2 c484 (.A0(net805),
    .A1(net260),
    .A2(net243),
    .A3(net145),
    .S0(clknet_1_1__leaf_net368),
    .S1(net699),
    .X(net380));
 sky130_fd_sc_hd__a2111oi_1 c485 (.A1(net219),
    .A2(net823),
    .B1(net257),
    .C1(net694),
    .D1(net991),
    .Y(net381));
 sky130_fd_sc_hd__sdfbbn_1 c486 (.CLK_N(clknet_4_12_0_clk),
    .D(net265),
    .RESET_B(net350),
    .SCD(net870),
    .SCE(clknet_1_0__leaf_net832),
    .SET_B(net927),
    .Q(net857));
 sky130_fd_sc_hd__sdfsbp_1 c487 (.CLK(clknet_4_12_0_clk),
    .D(net282),
    .SCD(net1005),
    .SCE(net273),
    .SET_B(net133),
    .Q(net383),
    .Q_N(net382));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net886),
    .A1(net383),
    .A2(net912),
    .A3(clknet_1_1__leaf_net849),
    .S0(clknet_1_0__leaf_net230),
    .S1(net685),
    .X(net384));
 sky130_fd_sc_hd__o2111ai_4 c489 (.A1(net841),
    .A2(net343),
    .B1(net838),
    .C1(net685),
    .D1(net847),
    .Y(net835));
 sky130_fd_sc_hd__mux4_4 c490 (.A0(net350),
    .A1(net370),
    .A2(net282),
    .A3(net145),
    .S0(net382),
    .S1(net835),
    .X(net385));
 sky130_fd_sc_hd__sdfstp_1 c491 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net368),
    .SCD(net383),
    .SCE(net935),
    .SET_B(net257),
    .Q(net386));
 sky130_fd_sc_hd__or4_1 c492 (.A(net670),
    .B(net847),
    .C(net840),
    .D(net700),
    .X(net853));
 sky130_fd_sc_hd__sdfbbp_1 c493 (.CLK(clknet_4_9_0_clk),
    .D(net145),
    .RESET_B(net1007),
    .SCD(net265),
    .SCE(net343),
    .SET_B(net931),
    .Q(net387));
 sky130_fd_sc_hd__and4bb_1 c494 (.A_N(net231),
    .B_N(net348),
    .C(net835),
    .D(net700),
    .X(net388));
 sky130_fd_sc_hd__a2111o_2 c495 (.A1(net910),
    .A2(net382),
    .B1(net386),
    .C1(net931),
    .D1(net701),
    .X(net389));
 sky130_fd_sc_hd__mux4_2 c496 (.A0(net356),
    .A1(net387),
    .A2(net389),
    .A3(net886),
    .S0(net281),
    .S1(net910),
    .X(net390));
 sky130_fd_sc_hd__mux4_2 c497 (.A0(net243),
    .A1(net264),
    .A2(net39),
    .A3(net834),
    .S0(net840),
    .S1(net699),
    .X(net391));
 sky130_fd_sc_hd__mux4_4 c498 (.A0(net26),
    .A1(net391),
    .A2(net21),
    .A3(net924),
    .S0(net887),
    .S1(net686),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net391),
    .A1(net386),
    .A2(net389),
    .A3(net885),
    .S0(net700),
    .S1(clknet_1_0__leaf_net702),
    .X(net393));
 sky130_fd_sc_hd__o2111ai_2 c500 (.A1(net389),
    .A2(net382),
    .B1(net929),
    .C1(net974),
    .D1(net704),
    .Y(net394));
 sky130_fd_sc_hd__a2111o_4 c501 (.A1(net394),
    .A2(net386),
    .B1(net311),
    .C1(net388),
    .D1(net700),
    .X(net395));
 sky130_fd_sc_hd__mux4_4 c502 (.A0(net386),
    .A1(net835),
    .A2(net273),
    .A3(net128),
    .S0(net858),
    .S1(net686),
    .X(net396));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net249),
    .A1(net835),
    .A2(net389),
    .A3(net821),
    .S0(net840),
    .S1(net705),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net311),
    .A1(net386),
    .A2(net397),
    .A3(net389),
    .S0(net877),
    .S1(net932),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net353),
    .A1(net388),
    .A2(net391),
    .A3(net26),
    .S0(net397),
    .S1(net707),
    .X(net399));
 sky130_fd_sc_hd__and2_1 c528 (.A(net66),
    .B(net306),
    .X(net400));
 sky130_fd_sc_hd__nor2b_4 c529 (.A(net74),
    .B_N(net297),
    .Y(net401));
 sky130_fd_sc_hd__nand2_4 c530 (.A(net188),
    .B(net64),
    .Y(net402));
 sky130_fd_sc_hd__nand2_4 c531 (.A(net933),
    .B(net306),
    .Y(net822));
 sky130_fd_sc_hd__or3b_2 c532 (.A(net306),
    .B(net763),
    .C_N(net402),
    .X(net403));
 sky130_fd_sc_hd__or2_1 c533 (.A(net79),
    .B(net822),
    .X(net404));
 sky130_fd_sc_hd__nand2_1 c534 (.A(net404),
    .B(net403),
    .Y(net405));
 sky130_fd_sc_hd__and2b_1 c535 (.A_N(net402),
    .B(net921),
    .X(net406));
 sky130_fd_sc_hd__nand4b_2 c536 (.A_N(net403),
    .B(net405),
    .C(net918),
    .D(net306),
    .Y(net407));
 sky130_fd_sc_hd__o2111a_2 c537 (.A1(net177),
    .A2(net306),
    .B1(net402),
    .C1(net292),
    .D1(net933),
    .X(net408));
 sky130_fd_sc_hd__and2b_1 c538 (.A_N(net406),
    .B(net404),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c539 (.A0(net407),
    .A1(net406),
    .A2(net403),
    .A3(net301),
    .S0(net400),
    .S1(net918),
    .X(net410));
 sky130_fd_sc_hd__and3b_1 c540 (.A_N(net301),
    .B(net402),
    .C(net407),
    .X(net411));
 sky130_fd_sc_hd__or4b_1 c541 (.A(net410),
    .B(net407),
    .C(net411),
    .D_N(net815),
    .X(net412));
 sky130_fd_sc_hd__mux4_2 c542 (.A0(net412),
    .A1(net406),
    .A2(net301),
    .A3(net75),
    .S0(net896),
    .S1(net64),
    .X(net413));
 sky130_fd_sc_hd__and4_4 c543 (.A(net405),
    .B(net406),
    .C(net413),
    .D(net75),
    .X(net833));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net400),
    .A1(net413),
    .A2(net408),
    .A3(net411),
    .S0(net833),
    .S1(net402),
    .X(net414));
 sky130_fd_sc_hd__nand4b_1 c545 (.A_N(net403),
    .B(net413),
    .C(net918),
    .D(net709),
    .Y(net415));
 sky130_fd_sc_hd__and3_1 c546 (.A(net921),
    .B(net411),
    .C(net407),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(net416),
    .A1(net298),
    .A2(net403),
    .A3(net833),
    .S0(net415),
    .S1(net413),
    .X(net417));
 sky130_fd_sc_hd__mux4_4 c548 (.A0(net415),
    .A1(net921),
    .A2(net412),
    .A3(net407),
    .S0(net402),
    .S1(net411),
    .X(net418));
 sky130_fd_sc_hd__nor4_1 c549 (.A(net413),
    .B(net411),
    .C(net410),
    .D(net667),
    .Y(net419));
 sky130_fd_sc_hd__and3b_1 c550 (.A_N(net322),
    .B(net185),
    .C(net676),
    .X(net420));
 sky130_fd_sc_hd__nand2_4 c551 (.A(net185),
    .B(net91),
    .Y(net421));
 sky130_fd_sc_hd__or2b_2 c552 (.A(net326),
    .B_N(net935),
    .X(net422));
 sky130_fd_sc_hd__and2_1 c553 (.A(net85),
    .B(net324),
    .X(net423));
 sky130_fd_sc_hd__nor3b_1 c554 (.A(net411),
    .B(net916),
    .C_N(net85),
    .Y(net424));
 sky130_fd_sc_hd__or3_2 c555 (.A(net423),
    .B(net420),
    .C(net919),
    .X(net425));
 sky130_fd_sc_hd__inv_16 c558_2 (.A(clknet_1_1__leaf_net673),
    .Y(net937));
 sky130_fd_sc_hd__buf_12 c557 (.A(clknet_1_0__leaf_net673),
    .X(net427));
 sky130_fd_sc_hd__clkinv_1 c316_7 (.A(net675),
    .Y(net942));
 sky130_fd_sc_hd__nor3b_4 c559 (.A(net217),
    .B(net896),
    .C_N(clknet_1_0__leaf_net427),
    .Y(net429));
 sky130_fd_sc_hd__mux4_4 c560 (.A0(net408),
    .A1(net941),
    .A2(net315),
    .A3(net195),
    .S0(clknet_1_0__leaf_net427),
    .S1(net671),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 c561 (.A(clknet_1_1__leaf_net758),
    .X(net431));
 sky130_fd_sc_hd__sdfbbn_1 c562 (.CLK_N(clknet_4_4_0_clk),
    .D(net296),
    .RESET_B(net421),
    .SCD(clknet_1_0__leaf_net427),
    .SCE(net422),
    .SET_B(net1000),
    .Q(net433),
    .Q_N(net432));
 sky130_fd_sc_hd__and3_2 c563 (.A(net940),
    .B(net774),
    .C(net677),
    .X(net434));
 sky130_fd_sc_hd__and3_4 c564 (.A(net425),
    .B(net423),
    .C(clknet_1_0__leaf_net434),
    .X(net435));
 sky130_fd_sc_hd__mux4_2 c565 (.A0(net342),
    .A1(clknet_1_0__leaf_net431),
    .A2(net422),
    .A3(net939),
    .S0(net898),
    .S1(net402),
    .X(net436));
 sky130_fd_sc_hd__nand4_4 c566 (.A(net421),
    .B(net238),
    .C(net679),
    .D(net931),
    .Y(net437));
 sky130_fd_sc_hd__nor4_4 c567 (.A(net437),
    .B(net408),
    .C(clknet_1_0__leaf_net434),
    .D(net676),
    .Y(net438));
 sky130_fd_sc_hd__sdfstp_1 c568 (.CLK(clknet_4_4_0_clk),
    .D(net430),
    .SCD(net425),
    .SCE(net437),
    .SET_B(clknet_1_0__leaf_net427),
    .Q(net439));
 sky130_fd_sc_hd__o2111ai_1 c569 (.A1(net315),
    .A2(clknet_1_0__leaf_net438),
    .B1(net439),
    .C1(net917),
    .D1(clknet_1_0__leaf_net427),
    .Y(net440));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net435),
    .A1(clknet_1_0__leaf_net438),
    .A2(net439),
    .A3(clknet_1_0__leaf_net434),
    .S0(net402),
    .S1(net327),
    .X(net441));
 sky130_fd_sc_hd__mux4_2 c571 (.A0(net439),
    .A1(net916),
    .A2(net423),
    .A3(net763),
    .S0(net408),
    .S1(net437),
    .X(net442));
 sky130_fd_sc_hd__or2b_1 c572 (.A(net201),
    .B_N(net0),
    .X(net443));
 sky130_fd_sc_hd__and4bb_4 c573 (.A_N(clknet_1_1__leaf_net232),
    .B_N(clknet_1_0__leaf_net431),
    .C(net298),
    .D(net822),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_4 c574 (.A(net625),
    .X(net444));
 sky130_fd_sc_hd__or3b_4 c575 (.A(net298),
    .B(clknet_1_0__leaf_net434),
    .C_N(net420),
    .X(net445));
 sky130_fd_sc_hd__inv_4 c576 (.A(net624),
    .Y(net446));
 sky130_fd_sc_hd__clkbuf_1 c577 (.A(net639),
    .X(net447));
 sky130_fd_sc_hd__or3_1 c578 (.A(net443),
    .B(net444),
    .C(clknet_1_0__leaf_net832),
    .X(net448));
 sky130_fd_sc_hd__o2111ai_4 c579 (.A1(net444),
    .A2(clknet_1_0__leaf_net427),
    .B1(net421),
    .C1(net915),
    .D1(net347),
    .Y(net449));
 sky130_fd_sc_hd__or3_4 c580 (.A(net446),
    .B(clknet_1_0__leaf_net445),
    .C(net964),
    .X(net450));
 sky130_fd_sc_hd__nor2_1 c581 (.A(clknet_1_1__leaf_net445),
    .B(net709),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 c582 (.A(net640),
    .Y(net452));
 sky130_fd_sc_hd__and3b_2 c583 (.A_N(net936),
    .B(clknet_1_0__leaf_net451),
    .C(net970),
    .X(net453));
 sky130_fd_sc_hd__nor3b_1 c584 (.A(net212),
    .B(clknet_1_0__leaf_net451),
    .C_N(net444),
    .Y(net454));
 sky130_fd_sc_hd__mux4_2 c585 (.A0(clknet_1_0__leaf_net454),
    .A1(clknet_1_1__leaf_net451),
    .A2(clknet_1_0__leaf_net434),
    .A3(net915),
    .S0(net324),
    .S1(clknet_1_0__leaf_net228),
    .X(net455));
 sky130_fd_sc_hd__nand3b_1 c586 (.A_N(clknet_1_1__leaf_net451),
    .B(clknet_1_1__leaf_net454),
    .C(clknet_1_0__leaf_net453),
    .Y(net456));
 sky130_fd_sc_hd__a2111oi_4 c587 (.A1(net452),
    .A2(net409),
    .B1(clknet_1_1__leaf_net451),
    .C1(clknet_1_0__leaf_net454),
    .D1(net446),
    .Y(net843));
 sky130_fd_sc_hd__and3b_4 c588 (.A_N(net449),
    .B(net444),
    .C(clknet_1_0__leaf_net843),
    .X(net457));
 sky130_fd_sc_hd__mux4_4 c589 (.A0(net946),
    .A1(clknet_1_0__leaf_net457),
    .A2(net452),
    .A3(clknet_1_0__leaf_net843),
    .S0(clknet_1_0__leaf_net454),
    .S1(net409),
    .X(net458));
 sky130_fd_sc_hd__mux4_4 c590 (.A0(net456),
    .A1(clknet_1_1__leaf_net454),
    .A2(net444),
    .A3(clknet_1_0__leaf_net457),
    .S0(clknet_1_0__leaf_net843),
    .S1(net710),
    .X(net459));
 sky130_fd_sc_hd__mux4_2 c591 (.A0(net447),
    .A1(clknet_1_1__leaf_net453),
    .A2(clknet_1_0__leaf_net457),
    .A3(clknet_1_1__leaf_net228),
    .S0(clknet_1_1__leaf_net454),
    .S1(net710),
    .X(net460));
 sky130_fd_sc_hd__a2111oi_2 c592 (.A1(net448),
    .A2(net821),
    .B1(clknet_1_0__leaf_net843),
    .C1(clknet_1_0__leaf_net454),
    .D1(net710),
    .Y(net461));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(clknet_1_0__leaf_net461),
    .A1(clknet_1_1__leaf_net457),
    .A2(net444),
    .A3(clknet_1_1__leaf_net454),
    .S0(net660),
    .S1(net665),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 c594 (.A(net756),
    .X(net463));
 sky130_fd_sc_hd__or3b_1 c595 (.A(net822),
    .B(net253),
    .C_N(net710),
    .X(net464));
 sky130_fd_sc_hd__or3b_1 c596 (.A(clknet_1_1__leaf_net431),
    .B(net463),
    .C_N(net23),
    .X(net465));
 sky130_fd_sc_hd__nor3_1 c597 (.A(net421),
    .B(net260),
    .C(net822),
    .Y(net466));
 sky130_fd_sc_hd__and4_4 c598 (.A(net788),
    .B(net21),
    .C(net348),
    .D(net969),
    .X(net467));
 sky130_fd_sc_hd__sdfbbn_1 c599 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net434),
    .RESET_B(net23),
    .SCD(net359),
    .SCE(net378),
    .SET_B(net920),
    .Q(net469),
    .Q_N(net468));
 sky130_fd_sc_hd__and3b_4 c600 (.A_N(net464),
    .B(clknet_1_0__leaf_net465),
    .C(net709),
    .X(net470));
 sky130_fd_sc_hd__or3_4 c601 (.A(clknet_1_0__leaf_net470),
    .B(net365),
    .C(net851),
    .X(net471));
 sky130_fd_sc_hd__o2111a_1 c602 (.A1(clknet_1_0__leaf_net471),
    .A2(net466),
    .B1(net467),
    .C1(clknet_1_0__leaf_net470),
    .D1(net890),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net361),
    .A1(clknet_1_0__leaf_net470),
    .A2(net833),
    .A3(clknet_1_0__leaf_net849),
    .S0(net464),
    .S1(net890),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net420),
    .A1(net359),
    .A2(clknet_1_0__leaf_net849),
    .A3(clknet_1_0__leaf_net470),
    .S0(clknet_1_0__leaf_net472),
    .S1(net711),
    .X(net474));
 sky130_fd_sc_hd__and4b_2 c605 (.A_N(net367),
    .B(clknet_1_1__leaf_net431),
    .C(net896),
    .D(clknet_1_0__leaf_net472),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net900),
    .A1(clknet_1_0__leaf_net471),
    .A2(clknet_1_0__leaf_net470),
    .A3(net444),
    .S0(net710),
    .S1(net711),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net366),
    .A1(net822),
    .A2(net378),
    .A3(net833),
    .S0(net889),
    .S1(clknet_1_1__leaf_net470),
    .X(net477));
 sky130_fd_sc_hd__sdfstp_1 c608 (.CLK(clknet_4_3_0_clk),
    .D(net476),
    .SCD(clknet_1_1__leaf_net472),
    .SCE(net972),
    .SET_B(net889),
    .Q(net478));
 sky130_fd_sc_hd__o2111ai_4 c609 (.A1(net807),
    .A2(net822),
    .B1(net890),
    .C1(net695),
    .D1(net712),
    .Y(net479));
 sky130_fd_sc_hd__mux4_2 c610 (.A0(net253),
    .A1(net478),
    .A2(net23),
    .A3(net479),
    .S0(clknet_1_1__leaf_net470),
    .S1(net712),
    .X(net480));
 sky130_fd_sc_hd__inv_2 c611 (.A(net756),
    .Y(net481));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net481),
    .A1(net788),
    .A2(net479),
    .A3(net833),
    .S0(clknet_1_0__leaf_net849),
    .S1(clknet_1_1__leaf_net674),
    .X(net482));
 sky130_fd_sc_hd__mux4_2 c613 (.A0(net455),
    .A1(net479),
    .A2(net900),
    .A3(clknet_1_0__leaf_net470),
    .S0(net712),
    .S1(net714),
    .X(net483));
 sky130_fd_sc_hd__mux4_4 c614 (.A0(net929),
    .A1(net479),
    .A2(clknet_1_1__leaf_net434),
    .A3(clknet_1_1__leaf_net471),
    .S0(clknet_1_0__leaf_net674),
    .S1(net713),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net327),
    .A1(clknet_1_1__leaf_net457),
    .A2(net479),
    .A3(clknet_1_0__leaf_net843),
    .S0(net361),
    .S1(net715),
    .X(net485));
 sky130_fd_sc_hd__o2111a_1 c616 (.A1(clknet_1_1__leaf_net843),
    .A2(net835),
    .B1(clknet_1_1__leaf_net849),
    .C1(net133),
    .D1(clknet_1_0__leaf_net703),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net348),
    .A1(net264),
    .A2(net915),
    .A3(net971),
    .S0(clknet_1_1__leaf_net843),
    .S1(net934),
    .X(net487));
 sky130_fd_sc_hd__sdfbbp_1 c618 (.CLK(clknet_4_12_0_clk),
    .D(net128),
    .RESET_B(net878),
    .SCD(net273),
    .SCE(net975),
    .SET_B(net706),
    .Q(net489),
    .Q_N(net488));
 sky130_fd_sc_hd__mux4_4 c619 (.A0(net257),
    .A1(net397),
    .A2(net128),
    .A3(net835),
    .S0(clknet_1_0__leaf_net824),
    .S1(clknet_1_0__leaf_net702),
    .X(net490));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net800),
    .A1(net802),
    .A2(net764),
    .A3(net3),
    .S0(net778),
    .S1(net798),
    .X(net0));
 sky130_fd_sc_hd__o2111a_1 c620 (.A1(net467),
    .A2(clknet_1_1__leaf_net427),
    .B1(net920),
    .C1(net658),
    .D1(net931),
    .X(net491));
 sky130_fd_sc_hd__a2111oi_0 c621 (.A1(clknet_1_1__leaf_net470),
    .A2(net91),
    .B1(net823),
    .C1(clknet_1_1__leaf_net427),
    .D1(net709),
    .Y(net492));
 sky130_fd_sc_hd__mux4_2 c622 (.A0(net912),
    .A1(net264),
    .A2(clknet_1_1__leaf_net427),
    .A3(net771),
    .S0(net665),
    .S1(net1000),
    .X(net493));
 sky130_fd_sc_hd__mux4_2 c623 (.A0(net491),
    .A1(net910),
    .A2(net934),
    .A3(net912),
    .S0(clknet_1_1__leaf_net427),
    .S1(net877),
    .X(net826));
 sky130_fd_sc_hd__mux4_4 c624 (.A0(net39),
    .A1(net489),
    .A2(net884),
    .A3(net21),
    .S0(net912),
    .S1(net706),
    .X(net494));
 sky130_fd_sc_hd__mux4_4 c625 (.A0(net912),
    .A1(net273),
    .A2(net133),
    .A3(net884),
    .S0(clknet_1_1__leaf_net702),
    .S1(net718),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net264),
    .A1(clknet_1_0__leaf_net487),
    .A2(net910),
    .A3(clknet_1_1__leaf_net470),
    .S0(net932),
    .S1(net718),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(clknet_1_0__leaf_net849),
    .A1(net833),
    .A2(clknet_1_1__leaf_net843),
    .A3(net264),
    .S0(net931),
    .S1(net716),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net784),
    .A1(clknet_1_0__leaf_net492),
    .A2(net920),
    .A3(net488),
    .S0(clknet_1_0__leaf_net720),
    .S1(clknet_1_0__leaf_net721),
    .X(net498));
 sky130_fd_sc_hd__mux4_4 c629 (.A0(net821),
    .A1(net273),
    .A2(clknet_1_1__leaf_net702),
    .A3(net718),
    .S0(clknet_1_1__leaf_net720),
    .S1(clknet_1_1__leaf_net721),
    .X(net499));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net787),
    .A1(net802),
    .A2(net798),
    .A3(net805),
    .S0(net808),
    .S1(net813),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net273),
    .A1(clknet_1_1__leaf_net492),
    .A2(net833),
    .A3(net284),
    .S0(net694),
    .S1(net722),
    .X(net500));
 sky130_fd_sc_hd__mux4_2 c631 (.A0(clknet_1_1__leaf_net427),
    .A1(clknet_1_1__leaf_net487),
    .A2(net784),
    .A3(net934),
    .S0(net719),
    .S1(clknet_1_0__leaf_net721),
    .X(net501));
 sky130_fd_sc_hd__mux4_4 c632 (.A0(net397),
    .A1(net932),
    .A2(clknet_1_1__leaf_net703),
    .A3(net708),
    .S0(net719),
    .S1(clknet_1_1__leaf_net721),
    .X(net502));
 sky130_fd_sc_hd__sdfbbn_1 c633 (.CLK_N(clknet_4_13_0_clk),
    .D(net915),
    .RESET_B(net493),
    .SCD(clknet_1_0__leaf_net487),
    .SCE(net929),
    .SET_B(net273),
    .Q(net503));
 sky130_fd_sc_hd__mux4_2 c634 (.A0(net503),
    .A1(net502),
    .A2(net39),
    .A3(clknet_1_0__leaf_net703),
    .S0(clknet_1_0__leaf_net720),
    .S1(clknet_1_1__leaf_net721),
    .X(net504));
 sky130_fd_sc_hd__mux4_2 c635 (.A0(net884),
    .A1(clknet_1_0__leaf_net492),
    .A2(net784),
    .A3(net257),
    .S0(net719),
    .S1(net726),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net498),
    .A1(net912),
    .A2(net854),
    .A3(net784),
    .S0(net724),
    .S1(net725),
    .X(net506));
 sky130_fd_sc_hd__mux4_4 c637 (.A0(net506),
    .A1(net884),
    .A2(clknet_1_1__leaf_net230),
    .A3(net699),
    .S0(net723),
    .S1(net727),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c64 (.A0(net801),
    .A1(net809),
    .A2(net802),
    .A3(net810),
    .S0(net811),
    .S1(net806),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net783),
    .A1(net775),
    .A2(net762),
    .A3(net779),
    .S0(net787),
    .S1(net820),
    .X(net3));
 sky130_fd_sc_hd__nor2_1 c66 (.A(net790),
    .B(net820),
    .Y(net4));
 sky130_fd_sc_hd__inv_6 c660 (.A(net628),
    .Y(net508));
 sky130_fd_sc_hd__nor2_1 c661 (.A(net190),
    .B(net763),
    .Y(net509));
 sky130_fd_sc_hd__buf_6 c662 (.A(net628),
    .X(net510));
 sky130_fd_sc_hd__or3b_1 c663 (.A(net510),
    .B(net509),
    .C_N(net667),
    .X(net511));
 sky130_fd_sc_hd__or2b_1 c664 (.A(net401),
    .B_N(net667),
    .X(net512));
 sky130_fd_sc_hd__or2b_2 c665 (.A(net815),
    .B_N(net667),
    .X(net513));
 sky130_fd_sc_hd__and3b_1 c666 (.A_N(net510),
    .B(net508),
    .C(net513),
    .X(net514));
 sky130_fd_sc_hd__and2b_1 c667 (.A_N(net509),
    .B(net508),
    .X(net515));
 sky130_fd_sc_hd__and3_2 c668 (.A(net292),
    .B(net510),
    .C(net512),
    .X(net516));
 sky130_fd_sc_hd__and2_1 c669 (.A(net515),
    .B(net513),
    .X(net517));
 sky130_fd_sc_hd__nor2b_2 c67 (.A(net771),
    .B_N(net780),
    .Y(net5));
 sky130_fd_sc_hd__nor3b_4 c670 (.A(net529),
    .B(net292),
    .C_N(net515),
    .Y(net518));
 sky130_fd_sc_hd__nor2b_1 c671 (.A(net517),
    .B_N(net516),
    .Y(net519));
 sky130_fd_sc_hd__mux4_1 c672 (.A0(net519),
    .A1(net514),
    .A2(net518),
    .A3(net529),
    .S0(net508),
    .S1(net510),
    .X(net520));
 sky130_fd_sc_hd__and3b_1 c673 (.A_N(net191),
    .B(net292),
    .C(net899),
    .X(net521));
 sky130_fd_sc_hd__or3_1 c674 (.A(net521),
    .B(net899),
    .C(net517),
    .X(net522));
 sky130_fd_sc_hd__mux4_2 c675 (.A0(net528),
    .A1(net191),
    .A2(net521),
    .A3(net529),
    .S0(net516),
    .S1(net510),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net1014),
    .A1(net518),
    .A2(net883),
    .A3(net896),
    .S0(net521),
    .S1(net996),
    .X(net524));
 sky130_fd_sc_hd__mux4_4 c677 (.A0(net519),
    .A1(net508),
    .A2(net518),
    .A3(net899),
    .S0(net523),
    .S1(net647),
    .X(net525));
 sky130_fd_sc_hd__nor3_1 c678 (.A(net523),
    .B(net519),
    .C(net646),
    .Y(net526));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net525),
    .A1(net522),
    .A2(net883),
    .A3(net899),
    .S0(net523),
    .S1(net646),
    .X(net527));
 sky130_fd_sc_hd__and2_1 c68 (.A(net5),
    .B(net935),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 c680 (.A(net647),
    .X(net528));
 sky130_fd_sc_hd__or2b_1 c681 (.A(net528),
    .B_N(net667),
    .X(net529));
 sky130_fd_sc_hd__nand3b_4 c682 (.A_N(net512),
    .B(net819),
    .C(net924),
    .Y(net530));
 sky130_fd_sc_hd__or3_2 c683 (.A(net522),
    .B(net514),
    .C(net401),
    .X(net531));
 sky130_fd_sc_hd__and3b_2 c684 (.A_N(net401),
    .B(net518),
    .C(net930),
    .X(net532));
 sky130_fd_sc_hd__nor3b_4 c685 (.A(net513),
    .B(net914),
    .C_N(net530),
    .Y(net533));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net514),
    .A1(net425),
    .A2(net512),
    .A3(net516),
    .S0(net815),
    .S1(net930),
    .X(net534));
 sky130_fd_sc_hd__and4_2 c687 (.A(net532),
    .B(net526),
    .C(net920),
    .D(net531),
    .X(net535));
 sky130_fd_sc_hd__o2111ai_1 c688 (.A1(net534),
    .A2(net425),
    .B1(net531),
    .C1(net516),
    .D1(net914),
    .Y(net536));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net526),
    .A1(net914),
    .A2(net532),
    .A3(net774),
    .S0(net899),
    .S1(net932),
    .X(net537));
 sky130_fd_sc_hd__and2b_1 c69 (.A_N(net5),
    .B(net808),
    .X(net7));
 sky130_fd_sc_hd__o2111a_1 c690 (.A1(net516),
    .A2(net401),
    .B1(net530),
    .C1(net649),
    .D1(net931),
    .X(net538));
 sky130_fd_sc_hd__nor4b_1 c691 (.A(net537),
    .B(net538),
    .C(net522),
    .D_N(net931),
    .Y(net539));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net914),
    .A1(net774),
    .A2(net538),
    .A3(net532),
    .S0(clknet_1_1__leaf_net438),
    .S1(net881),
    .X(net540));
 sky130_fd_sc_hd__mux4_4 c693 (.A0(net882),
    .A1(net526),
    .A2(net533),
    .A3(net535),
    .S0(net518),
    .S1(net679),
    .X(net541));
 sky130_fd_sc_hd__mux4_2 c694 (.A0(net402),
    .A1(net513),
    .A2(net195),
    .A3(net401),
    .S0(net518),
    .S1(net731),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net774),
    .A1(net532),
    .A2(net538),
    .A3(net649),
    .S0(net930),
    .S1(net731),
    .X(net543));
 sky130_fd_sc_hd__nor3b_1 c696 (.A(net543),
    .B(net195),
    .C_N(net935),
    .Y(net544));
 sky130_fd_sc_hd__mux4_2 c697 (.A0(net511),
    .A1(net938),
    .A2(net532),
    .A3(net195),
    .S0(net924),
    .S1(net731),
    .X(net545));
 sky130_fd_sc_hd__and4bb_1 c698 (.A_N(net511),
    .B_N(net829),
    .C(net401),
    .D(net731),
    .X(net546));
 sky130_fd_sc_hd__mux4_4 c699 (.A0(net544),
    .A1(net530),
    .A2(net535),
    .A3(clknet_1_1__leaf_net545),
    .S0(net542),
    .S1(net930),
    .X(net547));
 sky130_fd_sc_hd__and2_1 c70 (.A(net6),
    .B(net805),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(clknet_1_0__leaf_net545),
    .A1(net534),
    .A2(net530),
    .A3(net542),
    .S0(net932),
    .S1(net730),
    .X(net548));
 sky130_fd_sc_hd__nand4_4 c701 (.A(net442),
    .B(net402),
    .C(net542),
    .D(net930),
    .Y(net549));
 sky130_fd_sc_hd__a2111oi_1 c702 (.A1(net542),
    .A2(net546),
    .B1(net543),
    .C1(net899),
    .D1(net730),
    .Y(net550));
 sky130_fd_sc_hd__mux4_4 c703 (.A0(net550),
    .A1(clknet_1_1__leaf_net438),
    .A2(net549),
    .A3(net544),
    .S0(clknet_1_0__leaf_net547),
    .S1(net731),
    .X(net551));
 sky130_fd_sc_hd__mux4_2 c704 (.A0(clknet_1_0__leaf_net547),
    .A1(clknet_1_1__leaf_net230),
    .A2(net771),
    .A3(net195),
    .S0(net649),
    .S1(net732),
    .X(net552));
 sky130_fd_sc_hd__or4b_1 c705 (.A(net433),
    .B(net899),
    .C(net347),
    .D_N(net649),
    .X(net553));
 sky130_fd_sc_hd__or4b_2 c706 (.A(net937),
    .B(net531),
    .C(clknet_1_0__leaf_net547),
    .D_N(net930),
    .X(net554));
 sky130_fd_sc_hd__o2111a_2 c707 (.A1(net450),
    .A2(net532),
    .B1(net210),
    .C1(net666),
    .D1(net733),
    .X(net555));
 sky130_fd_sc_hd__sedfxbp_2 c708 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net440),
    .DE(net432),
    .SCD(net665),
    .SCE(net930),
    .Q(net557),
    .Q_N(net556));
 sky130_fd_sc_hd__o2111ai_4 c709 (.A1(net899),
    .A2(net917),
    .B1(net556),
    .C1(net649),
    .D1(net930),
    .Y(net558));
 sky130_fd_sc_hd__and2_0 c71 (.A(net803),
    .B(net815),
    .X(net9));
 sky130_fd_sc_hd__a2111o_2 c710 (.A1(net531),
    .A2(net780),
    .B1(net899),
    .C1(clknet_1_1__leaf_net440),
    .D1(net735),
    .X(net559));
 sky130_fd_sc_hd__or3_2 c711 (.A(net195),
    .B(net557),
    .C(net348),
    .X(net560));
 sky130_fd_sc_hd__sdfbbn_1 c712 (.CLK_N(clknet_4_5_0_clk),
    .D(net555),
    .RESET_B(net920),
    .SCD(net556),
    .SCE(net532),
    .SET_B(net1002),
    .Q(net561));
 sky130_fd_sc_hd__a2111oi_1 c713 (.A1(net535),
    .A2(clknet_1_1__leaf_net230),
    .B1(net899),
    .C1(net930),
    .D1(net734),
    .Y(net562));
 sky130_fd_sc_hd__sedfxbp_1 c714 (.CLK(clknet_4_6_0_clk),
    .D(net557),
    .DE(clknet_1_0__leaf_net824),
    .SCD(net324),
    .SCE(net347),
    .Q(net563));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net1013),
    .A1(net433),
    .A2(net195),
    .A3(net549),
    .S0(net556),
    .S1(net711),
    .X(net564));
 sky130_fd_sc_hd__sdfbbp_1 c716 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net461),
    .RESET_B(net532),
    .SCD(net1012),
    .SCE(net0),
    .SET_B(net771),
    .Q(net566),
    .Q_N(net565));
 sky130_fd_sc_hd__mux4_2 c717 (.A0(net896),
    .A1(net973),
    .A2(clknet_1_0__leaf_net562),
    .A3(net520),
    .S0(net734),
    .S1(net736),
    .X(net567));
 sky130_fd_sc_hd__a2111oi_4 c718 (.A1(net553),
    .A2(net432),
    .B1(net784),
    .C1(net566),
    .D1(net736),
    .Y(net568));
 sky130_fd_sc_hd__mux4_4 c719 (.A0(net558),
    .A1(net897),
    .A2(clknet_1_1__leaf_net547),
    .A3(net930),
    .S0(net736),
    .S1(net737),
    .X(net569));
 sky130_fd_sc_hd__and3b_2 c72 (.A_N(net784),
    .B(net8),
    .C(net787),
    .X(net838));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net771),
    .A1(net897),
    .A2(net556),
    .A3(net565),
    .S0(net729),
    .S1(net735),
    .X(net570));
 sky130_fd_sc_hd__o2111a_1 c721 (.A1(net570),
    .A2(net557),
    .B1(net774),
    .C1(net530),
    .D1(net738),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net570),
    .A1(clknet_1_1__leaf_net562),
    .A2(clknet_1_1__leaf_net547),
    .A3(net535),
    .S0(net897),
    .S1(net565),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net774),
    .A1(net568),
    .A2(net565),
    .A3(net711),
    .S0(net736),
    .S1(clknet_1_0__leaf_net739),
    .X(net573));
 sky130_fd_sc_hd__o2111a_4 c724 (.A1(net210),
    .A2(net558),
    .B1(net535),
    .C1(net560),
    .D1(clknet_1_1__leaf_net739),
    .X(net574));
 sky130_fd_sc_hd__sdfbbn_1 c725 (.CLK_N(clknet_4_5_0_clk),
    .D(net997),
    .RESET_B(clknet_1_0__leaf_net574),
    .SCD(net566),
    .SCE(net666),
    .SET_B(net736),
    .Q(net576),
    .Q_N(net575));
 sky130_fd_sc_hd__mux4_2 c726 (.A0(clknet_1_0__leaf_net465),
    .A1(net444),
    .A2(net467),
    .A3(net362),
    .S0(net829),
    .S1(net711),
    .X(net577));
 sky130_fd_sc_hd__a2111oi_1 c727 (.A1(net571),
    .A2(net566),
    .B1(net807),
    .C1(net560),
    .D1(net655),
    .Y(net578));
 sky130_fd_sc_hd__mux4_2 c728 (.A0(clknet_1_0__leaf_net429),
    .A1(net890),
    .A2(net812),
    .A3(net771),
    .S0(net549),
    .S1(net730),
    .X(net579));
 sky130_fd_sc_hd__mux4_4 c729 (.A0(net479),
    .A1(clknet_1_1__leaf_net574),
    .A2(net347),
    .A3(net890),
    .S0(net972),
    .S1(net711),
    .X(net580));
 sky130_fd_sc_hd__nor3b_2 c73 (.A(net817),
    .B(net7),
    .C_N(net925),
    .Y(net10));
 sky130_fd_sc_hd__mux4_2 c730 (.A0(clknet_1_1__leaf_net429),
    .A1(net348),
    .A2(net546),
    .A3(net309),
    .S0(net933),
    .S1(net711),
    .X(net581));
 sky130_fd_sc_hd__a2111o_1 c731 (.A1(net566),
    .A2(net804),
    .B1(net347),
    .C1(clknet_1_1__leaf_net465),
    .D1(clknet_1_1__leaf_net740),
    .X(net582));
 sky130_fd_sc_hd__a2111o_2 c732 (.A1(clknet_1_1__leaf_net547),
    .A2(net924),
    .B1(net565),
    .C1(net735),
    .D1(clknet_1_0__leaf_net741),
    .X(net583));
 sky130_fd_sc_hd__a2111oi_1 c733 (.A1(net573),
    .A2(net379),
    .B1(net467),
    .C1(net736),
    .D1(clknet_1_0__leaf_net740),
    .Y(net584));
 sky130_fd_sc_hd__a2111o_4 c734 (.A1(net530),
    .A2(net890),
    .B1(clknet_1_1__leaf_net429),
    .C1(net767),
    .D1(net880),
    .X(net585));
 sky130_fd_sc_hd__mux4_4 c735 (.A0(net379),
    .A1(net348),
    .A2(net568),
    .A3(net890),
    .S0(clknet_1_1__leaf_net429),
    .S1(net711),
    .X(net586));
 sky130_fd_sc_hd__sdfbbn_1 c736 (.CLK_N(clknet_4_7_0_clk),
    .D(net1004),
    .RESET_B(net549),
    .SCD(clknet_1_1__leaf_net824),
    .SCE(net920),
    .SET_B(net736),
    .Q(net588),
    .Q_N(net587));
 sky130_fd_sc_hd__o2111a_1 c737 (.A1(net575),
    .A2(net379),
    .B1(net763),
    .C1(net657),
    .D1(clknet_1_0__leaf_net741),
    .X(net589));
 sky130_fd_sc_hd__sdfbbp_1 c738 (.CLK(clknet_4_7_0_clk),
    .D(net530),
    .RESET_B(net444),
    .SCD(clknet_1_1__leaf_net586),
    .SCE(net657),
    .SET_B(clknet_1_1__leaf_net741),
    .Q(net590));
 sky130_fd_sc_hd__mux4_4 c739 (.A0(net560),
    .A1(net589),
    .A2(net920),
    .A3(net890),
    .S0(clknet_1_1__leaf_net230),
    .S1(clknet_1_0__leaf_net577),
    .X(net591));
 sky130_fd_sc_hd__and4bb_1 c74 (.A_N(net2),
    .B_N(net6),
    .C(net10),
    .D(net925),
    .X(net11));
 sky130_fd_sc_hd__sdfbbn_2 c740 (.CLK_N(clknet_4_6_0_clk),
    .D(net546),
    .RESET_B(net1017),
    .SCD(net0),
    .SCE(net924),
    .SET_B(net998),
    .Q(net593),
    .Q_N(net592));
 sky130_fd_sc_hd__sdfbbn_1 c741 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net586),
    .RESET_B(net557),
    .SCD(net593),
    .SCE(net890),
    .SET_B(net998),
    .Q(net595),
    .Q_N(net594));
 sky130_fd_sc_hd__a2111oi_0 c742 (.A1(net584),
    .A2(net21),
    .B1(net594),
    .C1(net592),
    .D1(net742),
    .Y(net596));
 sky130_fd_sc_hd__mux4_4 c743 (.A0(net595),
    .A1(net780),
    .A2(net378),
    .A3(net592),
    .S0(net730),
    .S1(net736),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net362),
    .A1(net590),
    .A2(net587),
    .A3(net593),
    .S0(net594),
    .S1(clknet_1_1__leaf_net596),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net568),
    .A1(net581),
    .A2(net530),
    .A3(clknet_1_1__leaf_net596),
    .S0(net595),
    .S1(net592),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net324),
    .A1(net597),
    .A2(net593),
    .A3(net566),
    .S0(net594),
    .S1(net744),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_1__leaf_net577),
    .A1(net595),
    .A2(net444),
    .A3(net592),
    .S0(net600),
    .S1(net743),
    .X(net601));
 sky130_fd_sc_hd__mux4_4 c748 (.A0(net588),
    .A1(clknet_1_0__leaf_net582),
    .A2(net469),
    .A3(net533),
    .S0(net829),
    .S1(net745),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(clknet_1_1__leaf_net230),
    .A1(net260),
    .A2(net812),
    .A3(net533),
    .S0(net784),
    .S1(clknet_1_0__leaf_net596),
    .X(net603));
 sky130_fd_sc_hd__nor3_2 c75 (.A(net7),
    .B(net4),
    .C(net925),
    .Y(net12));
 sky130_fd_sc_hd__mux4_4 c750 (.A0(net533),
    .A1(net260),
    .A2(clknet_1_1__leaf_net824),
    .A3(net347),
    .S0(net727),
    .S1(net746),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net602),
    .A1(clknet_1_0__leaf_net596),
    .A2(clknet_1_1__leaf_net230),
    .A3(net717),
    .S0(net728),
    .S1(net747),
    .X(net605));
 sky130_fd_sc_hd__mux4_4 c752 (.A0(net593),
    .A1(net829),
    .A2(net468),
    .A3(net932),
    .S0(net748),
    .S1(net749),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net469),
    .A1(net606),
    .A2(net260),
    .A3(net924),
    .S0(net467),
    .S1(net728),
    .X(net607));
 sky130_fd_sc_hd__mux4_2 c754 (.A0(net133),
    .A1(net21),
    .A2(clknet_1_0__leaf_net824),
    .A3(net717),
    .S0(net728),
    .S1(net747),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net549),
    .A1(net600),
    .A2(net593),
    .A3(net855),
    .S0(net763),
    .S1(net1010),
    .X(net609));
 sky130_fd_sc_hd__mux4_4 c756 (.A0(clknet_1_0__leaf_net824),
    .A1(net661),
    .A2(net706),
    .A3(net726),
    .S0(net728),
    .S1(net747),
    .X(net610));
 sky130_fd_sc_hd__mux4_4 c757 (.A0(clknet_1_1__leaf_net582),
    .A1(net133),
    .A2(net592),
    .A3(net932),
    .S0(net707),
    .S1(net747),
    .X(net611));
 sky130_fd_sc_hd__mux4_2 c758 (.A0(net607),
    .A1(clknet_1_0__leaf_net611),
    .A2(net549),
    .A3(net920),
    .S0(clknet_1_1__leaf_net824),
    .S1(net747),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net593),
    .A1(net717),
    .A2(net725),
    .A3(net727),
    .S0(net749),
    .S1(net750),
    .X(net613));
 sky130_fd_sc_hd__nand3b_1 c76 (.A_N(net780),
    .B(net803),
    .C(net925),
    .Y(net13));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net533),
    .A1(net971),
    .A2(net613),
    .A3(net696),
    .S0(net747),
    .S1(net753),
    .X(net614));
 sky130_fd_sc_hd__mux4_4 c761 (.A0(net613),
    .A1(clknet_1_1__leaf_net611),
    .A2(net707),
    .A3(net727),
    .S0(net733),
    .S1(net747),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net0),
    .A1(net467),
    .A2(net614),
    .A3(clknet_1_0__leaf_net824),
    .S0(net855),
    .S1(net750),
    .X(net616));
 sky130_fd_sc_hd__mux4_4 c763 (.A0(net467),
    .A1(net613),
    .A2(net747),
    .A3(net748),
    .S0(net752),
    .S1(net754),
    .X(net617));
 sky130_fd_sc_hd__mux4_4 c764 (.A0(net615),
    .A1(net617),
    .A2(net614),
    .A3(clknet_1_0__leaf_net824),
    .S0(net728),
    .S1(net751),
    .X(net618));
 sky130_fd_sc_hd__or2_2 c77 (.A(net9),
    .B(net11),
    .X(net14));
 sky130_fd_sc_hd__nand3_2 c78 (.A(net808),
    .B(net13),
    .C(net925),
    .Y(net15));
 sky130_fd_sc_hd__and2_4 c79 (.A(net9),
    .B(net4),
    .X(net16));
 sky130_fd_sc_hd__and4b_4 c80 (.A_N(net12),
    .B(net14),
    .C(net16),
    .D(net925),
    .X(net17));
 sky130_fd_sc_hd__mux4_2 c81 (.A0(net6),
    .A1(net13),
    .A2(net10),
    .A3(net11),
    .S0(net817),
    .S1(net5),
    .X(net18));
 sky130_fd_sc_hd__nor3b_1 c82 (.A(net16),
    .B(net3),
    .C_N(net925),
    .Y(net19));
 sky130_fd_sc_hd__nand2b_2 c83 (.A_N(net13),
    .B(net14),
    .Y(net20));
 sky130_fd_sc_hd__mux4_2 c84 (.A0(net4),
    .A1(net11),
    .A2(net15),
    .A3(net775),
    .S0(net925),
    .S1(net20),
    .X(net21));
 sky130_fd_sc_hd__a2111oi_4 c85 (.A1(net8),
    .A2(net925),
    .B1(net18),
    .C1(net2),
    .D1(net20),
    .Y(net22));
 sky130_fd_sc_hd__mux4_2 c86 (.A0(net21),
    .A1(net6),
    .A2(net15),
    .A3(net20),
    .S0(net16),
    .S1(net923),
    .X(net23));
 sky130_fd_sc_hd__a2111o_4 c87 (.A1(net22),
    .A2(net20),
    .B1(net16),
    .C1(net17),
    .D1(net820),
    .X(net24));
 sky130_fd_sc_hd__and2_1 c88 (.A(net8),
    .B(net19),
    .X(net25));
 sky130_fd_sc_hd__and2_2 c89 (.A(net10),
    .B(net19),
    .X(net26));
 sky130_fd_sc_hd__nor2_1 c90 (.A(net776),
    .B(net25),
    .Y(net27));
 sky130_fd_sc_hd__and2_2 c91 (.A(net811),
    .B(net27),
    .X(net28));
 sky130_fd_sc_hd__nor2_1 c92 (.A(net27),
    .B(net25),
    .Y(net29));
 sky130_fd_sc_hd__and2_1 c93 (.A(net25),
    .B(net810),
    .X(net30));
 sky130_fd_sc_hd__nand2b_4 c94 (.A_N(net790),
    .B(net28),
    .Y(net31));
 sky130_fd_sc_hd__or3_4 c95 (.A(net19),
    .B(net24),
    .C(net31),
    .X(net32));
 sky130_fd_sc_hd__o2111a_1 c96 (.A1(net30),
    .A2(net20),
    .B1(net19),
    .C1(net32),
    .D1(net31),
    .X(net33));
 sky130_fd_sc_hd__nor2_1 c97 (.A(net29),
    .B(net32),
    .Y(net34));
 sky130_fd_sc_hd__or4b_4 c98 (.A(net34),
    .B(net33),
    .C(net32),
    .D_N(net28),
    .X(net869));
 sky130_fd_sc_hd__nand3_1 c99 (.A(net810),
    .B(net28),
    .C(net32),
    .Y(net35));
 sky130_fd_sc_hd__or4_1 merge765 (.A(net422),
    .B(net322),
    .C(net420),
    .D(net667),
    .X(net619));
 sky130_fd_sc_hd__sedfxtp_1 merge766 (.CLK(clknet_4_10_0_clk),
    .D(net56),
    .DE(net48),
    .SCD(net872),
    .SCE(net680),
    .Q(net620));
 sky130_fd_sc_hd__sedfxtp_4 merge767 (.CLK(clknet_4_1_0_clk),
    .D(net224),
    .DE(net774),
    .SCD(clknet_1_1__leaf_net341),
    .SCE(clknet_1_0__leaf_net345),
    .Q(net621));
 sky130_fd_sc_hd__mux4_1 merge768 (.A0(net239),
    .A1(net923),
    .A2(net252),
    .A3(net128),
    .S0(net247),
    .S1(net682),
    .X(net622));
 sky130_fd_sc_hd__mux4_2 merge769 (.A0(clknet_1_0__leaf_net429),
    .A1(clknet_1_1__leaf_net457),
    .A2(clknet_1_1__leaf_net832),
    .A3(net479),
    .S0(net296),
    .S1(net654),
    .X(net623));
 sky130_fd_sc_hd__sdfbbp_1 merge770 (.CLK(clknet_4_1_0_clk),
    .D(net917),
    .RESET_B(net833),
    .SCD(net965),
    .SCE(net807),
    .SET_B(net659),
    .Q(net625),
    .Q_N(net624));
 sky130_fd_sc_hd__nand4b_1 merge771 (.A_N(net124),
    .B(net845),
    .C(net83),
    .D(net112),
    .Y(net626));
 sky130_fd_sc_hd__or4b_1 merge772 (.A(net184),
    .B(net311),
    .C(net317),
    .D_N(net319),
    .X(net627));
 sky130_fd_sc_hd__inv_4 merge773 (.A(net647),
    .Y(net628));
 sky130_fd_sc_hd__sdfbbn_2 merge774 (.CLK_N(clknet_4_12_0_clk),
    .D(net316),
    .RESET_B(net21),
    .SCD(net219),
    .SCE(net889),
    .SET_B(net644),
    .Q(net630),
    .Q_N(net629));
 sky130_fd_sc_hd__nand4b_1 merge775 (.A_N(net809),
    .B(net888),
    .C(net221),
    .D(net201),
    .Y(net631));
 sky130_fd_sc_hd__sdfbbn_1 merge776 (.CLK_N(clknet_4_0_0_clk),
    .D(net121),
    .RESET_B(net776),
    .SCD(net69),
    .SCE(net891),
    .SET_B(net137),
    .Q(net633),
    .Q_N(net632));
 sky130_fd_sc_hd__sdfbbp_1 merge777 (.CLK(clknet_4_8_0_clk),
    .D(net47),
    .RESET_B(net24),
    .SCD(net155),
    .SCE(net866),
    .SET_B(net992),
    .Q(net635),
    .Q_N(net634));
 sky130_fd_sc_hd__mux4_1 merge778 (.A0(net77),
    .A1(clknet_1_0__leaf_net849),
    .A2(net915),
    .A3(net989),
    .S0(net208),
    .S1(net888),
    .X(net636));
 sky130_fd_sc_hd__o2111a_1 merge779 (.A1(net1016),
    .A2(net209),
    .B1(net222),
    .C1(clknet_1_0__leaf_net233),
    .D1(net206),
    .X(net637));
 sky130_fd_sc_hd__mux4_4 merge780 (.A0(net942),
    .A1(clknet_1_0__leaf_net230),
    .A2(net219),
    .A3(clknet_1_0__leaf_net339),
    .S0(net340),
    .S1(net904),
    .X(net638));
 sky130_fd_sc_hd__sdfbbn_1 merge781 (.CLK_N(clknet_4_1_0_clk),
    .D(net409),
    .RESET_B(clknet_1_0__leaf_net824),
    .SCD(clknet_1_0__leaf_net451),
    .SCE(clknet_1_0__leaf_net228),
    .SET_B(net64),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net408),
    .A1(net422),
    .A2(clknet_1_0__leaf_net427),
    .A3(net902),
    .S0(net186),
    .S1(net317),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(clknet_1_1__leaf_net345),
    .A1(net945),
    .A2(net915),
    .A3(net424),
    .S0(net422),
    .S1(net931),
    .X(net642));
 sky130_fd_sc_hd__nor4_1 merge784 (.A(net75),
    .B(net419),
    .C(net401),
    .D(net819),
    .Y(net643));
 sky130_fd_sc_hd__dfrbp_1 merge785 (.CLK(clknet_4_9_0_clk),
    .D(net256),
    .RESET_B(net261),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__dfrbp_2 merge786 (.CLK(clknet_4_4_0_clk),
    .D(net643),
    .RESET_B(net524),
    .Q(net647),
    .Q_N(net646));
 sky130_fd_sc_hd__dfrtn_1 merge787 (.CLK_N(clknet_4_9_0_clk),
    .D(net380),
    .RESET_B(net381),
    .Q(net858));
 sky130_fd_sc_hd__nand2b_1 merge788 (.A_N(net436),
    .B(net441),
    .Y(net648));
 sky130_fd_sc_hd__dfrtp_4 merge789 (.CLK(clknet_4_5_0_clk),
    .D(net536),
    .RESET_B(net548),
    .Q(net649));
 sky130_fd_sc_hd__dfrtp_1 merge790 (.CLK(clknet_4_11_0_clk),
    .RESET_B(net288),
    .Q(net290));
 sky130_fd_sc_hd__and2_1 merge791 (.A(net331),
    .B(net332),
    .X(net650));
 sky130_fd_sc_hd__dfrtp_1 merge792 (.CLK(clknet_4_8_0_clk),
    .D(net156),
    .RESET_B(net157),
    .Q(net651));
 sky130_fd_sc_hd__dfsbp_1 merge793 (.CLK(clknet_4_2_0_clk),
    .D(net139),
    .SET_B(net142),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__dfsbp_1 merge794 (.CLK(clknet_4_6_0_clk),
    .D(net473),
    .SET_B(net474),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__dfstp_1 merge795 (.CLK(clknet_4_2_0_clk),
    .D(net352),
    .Q(net355));
 sky130_fd_sc_hd__dfstp_2 merge796 (.CLK(clknet_4_3_0_clk),
    .D(net371),
    .SET_B(net364),
    .Q(net851));
 sky130_fd_sc_hd__dfstp_1 merge797 (.CLK(clknet_4_7_0_clk),
    .D(net583),
    .SET_B(net585),
    .Q(net657));
 sky130_fd_sc_hd__dlrbn_1 merge798 (.D(net486),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net490),
    .Q(net658));
 sky130_fd_sc_hd__dlrbn_1 merge799 (.D(net122),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net123),
    .Q_N(net659));
 sky130_fd_sc_hd__dlrbp_1 merge800 (.D(net618),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net609),
    .Q(net661));
 sky130_fd_sc_hd__dlrbp_2 merge801 (.D(net237),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net631),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__dlrtn_1 merge802 (.D(net57),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net60),
    .Q(net664));
 sky130_fd_sc_hd__dlrtn_2 merge803 (.D(net459),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net460),
    .Q(net665));
 sky130_fd_sc_hd__dlrtn_1 merge804 (.D(net554),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net559),
    .Q(net666));
 sky130_fd_sc_hd__dlrtp_1 merge805 (.D(net417),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net418),
    .Q(net667));
 sky130_fd_sc_hd__dlrtp_1 merge806 (.D(net274),
    .GATE(clknet_4_11_0_clk),
    .Q(net286));
 sky130_fd_sc_hd__dlrtp_1 merge807 (.D(net172),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net173),
    .Q(net669));
 sky130_fd_sc_hd__edfxbp_1 merge808 (.CLK(clknet_4_1_0_clk),
    .D(net333),
    .Q(net334),
    .Q_N(net670));
 sky130_fd_sc_hd__edfxtp_1 merge809 (.CLK(clknet_4_0_0_clk),
    .D(net140),
    .DE(net626),
    .Q(net672));
 sky130_fd_sc_hd__sdlclkp_1 merge810 (.CLK(clknet_4_1_0_clk),
    .GATE(net619),
    .SCE(net641),
    .GCLK(net673));
 sky130_fd_sc_hd__sdlclkp_2 merge811 (.CLK(clknet_4_6_0_clk),
    .GATE(net483),
    .SCE(net475),
    .GCLK(net674));
 sky130_fd_sc_hd__sdlclkp_4 merge812 (.CLK(clknet_4_0_0_clk),
    .GATE(net637),
    .SCE(net638),
    .GCLK(net675));
 sky130_fd_sc_hd__dfrbp_1 merge813 (.CLK(clknet_4_1_0_clk),
    .D(net627),
    .RESET_B(net325),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dfrbp_1 merge814 (.CLK(clknet_4_11_0_clk),
    .D(net395),
    .RESET_B(net175),
    .Q(net836),
    .Q_N(net678));
 sky130_fd_sc_hd__dfrtn_1 merge815 (.CLK_N(clknet_4_1_0_clk),
    .D(net648),
    .RESET_B(net650),
    .Q(net679));
 sky130_fd_sc_hd__dfxbp_1 s816 (.CLK(clknet_4_10_0_clk),
    .D(net58),
    .Q(net681),
    .Q_N(net680));
 sky130_fd_sc_hd__dfxbp_1 s817 (.CLK(clknet_4_8_0_clk),
    .D(net141),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__dfxtp_1 s818 (.CLK(clknet_4_10_0_clk),
    .D(net159),
    .Q(net684));
 sky130_fd_sc_hd__dfxtp_2 s819 (.CLK(clknet_4_8_0_clk),
    .D(net161),
    .Q(net685));
 sky130_fd_sc_hd__dfxtp_1 s820 (.CLK(clknet_4_8_0_clk),
    .D(net163),
    .Q(net686));
 sky130_fd_sc_hd__dlclkp_1 s821 (.CLK(clknet_4_10_0_clk),
    .GATE(net164),
    .GCLK(net687));
 sky130_fd_sc_hd__dlclkp_2 s822 (.CLK(clknet_4_10_0_clk),
    .GATE(net174),
    .GCLK(net688));
 sky130_fd_sc_hd__dlclkp_4 s823 (.CLK(clknet_4_10_0_clk),
    .GATE(net176),
    .GCLK(net689));
 sky130_fd_sc_hd__dlxbn_1 s824 (.D(net234),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net691),
    .Q_N(net690));
 sky130_fd_sc_hd__dlxbn_1 s825 (.D(net236),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net693),
    .Q_N(net692));
 sky130_fd_sc_hd__dlxbp_1 s826 (.D(net241),
    .GATE(clknet_4_2_0_clk),
    .Q(net877),
    .Q_N(net694));
 sky130_fd_sc_hd__dlxtn_1 s827 (.D(net244),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net856));
 sky130_fd_sc_hd__dlxtn_1 s828 (.D(net280),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net850));
 sky130_fd_sc_hd__dlxtn_2 s829 (.D(net285),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net847));
 sky130_fd_sc_hd__dlxtp_1 s830 (.D(net287),
    .GATE(clknet_4_9_0_clk),
    .Q(net840));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s831 (.D(net289),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net876));
 sky130_fd_sc_hd__dfxbp_2 s832 (.CLK(clknet_4_0_0_clk),
    .D(net328),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__dfxbp_1 s833 (.CLK(clknet_4_0_0_clk),
    .D(net329),
    .Q(net698),
    .Q_N(net697));
 sky130_fd_sc_hd__dfxtp_1 s834 (.CLK(clknet_4_9_0_clk),
    .D(net377),
    .Q(net699));
 sky130_fd_sc_hd__dfxtp_1 s835 (.CLK(clknet_4_11_0_clk),
    .D(net384),
    .Q(net700));
 sky130_fd_sc_hd__dfxtp_1 s836 (.CLK(clknet_4_12_0_clk),
    .D(net385),
    .Q(net701));
 sky130_fd_sc_hd__dlclkp_1 s837 (.CLK(clknet_4_11_0_clk),
    .GATE(net390),
    .GCLK(net702));
 sky130_fd_sc_hd__dlclkp_2 s838 (.CLK(clknet_4_12_0_clk),
    .GATE(net392),
    .GCLK(net703));
 sky130_fd_sc_hd__dlclkp_4 s839 (.CLK(clknet_4_11_0_clk),
    .GATE(net393),
    .GCLK(net704));
 sky130_fd_sc_hd__dlxbn_1 s840 (.D(net396),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net705));
 sky130_fd_sc_hd__dlxbn_1 s841 (.D(net398),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dlxbp_1 s842 (.D(net399),
    .GATE(clknet_4_14_0_clk),
    .Q(net879),
    .Q_N(net708));
 sky130_fd_sc_hd__dlxtn_2 s843 (.D(net414),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net709));
 sky130_fd_sc_hd__dlxtn_1 s844 (.D(net458),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net710));
 sky130_fd_sc_hd__dlxtn_4 s845 (.D(net462),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net711));
 sky130_fd_sc_hd__dlxtp_1 s846 (.D(net477),
    .GATE(clknet_4_3_0_clk),
    .Q(net712));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s847 (.D(net480),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net713));
 sky130_fd_sc_hd__dfxbp_1 s848 (.CLK(clknet_4_6_0_clk),
    .D(net482),
    .Q(net714));
 sky130_fd_sc_hd__dfxbp_1 s849 (.CLK(clknet_4_6_0_clk),
    .D(net484),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__dfxtp_1 s850 (.CLK(clknet_4_13_0_clk),
    .D(net485),
    .Q(net717));
 sky130_fd_sc_hd__dfxtp_1 s851 (.CLK(clknet_4_12_0_clk),
    .D(net494),
    .Q(net718));
 sky130_fd_sc_hd__dfxtp_1 s852 (.CLK(clknet_4_14_0_clk),
    .D(net495),
    .Q(net719));
 sky130_fd_sc_hd__dlclkp_1 s853 (.CLK(clknet_4_12_0_clk),
    .GATE(net496),
    .GCLK(net720));
 sky130_fd_sc_hd__dlclkp_2 s854 (.CLK(clknet_4_13_0_clk),
    .GATE(net497),
    .GCLK(net721));
 sky130_fd_sc_hd__dlclkp_4 s855 (.CLK(clknet_4_14_0_clk),
    .GATE(net499),
    .GCLK(net722));
 sky130_fd_sc_hd__dlxbn_1 s856 (.D(net500),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net723));
 sky130_fd_sc_hd__dlxbn_1 s857 (.D(net501),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net724));
 sky130_fd_sc_hd__dlxbp_1 s858 (.D(net504),
    .GATE(clknet_4_15_0_clk),
    .Q(net726),
    .Q_N(net725));
 sky130_fd_sc_hd__dlxtn_1 s859 (.D(net505),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net727));
 sky130_fd_sc_hd__dlxtn_2 s860 (.D(net507),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net728));
 sky130_fd_sc_hd__dlxtn_1 s861 (.D(net527),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net729));
 sky130_fd_sc_hd__dlxtp_1 s862 (.D(net540),
    .GATE(clknet_4_5_0_clk),
    .Q(net730));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s863 (.D(net541),
    .SLEEP_B(clknet_4_4_0_clk),
    .Q(net731));
 sky130_fd_sc_hd__dfxbp_1 s864 (.CLK(clknet_4_5_0_clk),
    .D(net551),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__dfxbp_1 s865 (.CLK(clknet_4_5_0_clk),
    .D(net552),
    .Q(net735),
    .Q_N(net734));
 sky130_fd_sc_hd__dfxtp_4 s866 (.CLK(clknet_4_6_0_clk),
    .D(net564),
    .Q(net736));
 sky130_fd_sc_hd__dfxtp_1 s867 (.CLK(clknet_4_5_0_clk),
    .D(net567),
    .Q(net737));
 sky130_fd_sc_hd__dfxtp_1 s868 (.CLK(clknet_4_5_0_clk),
    .D(net569),
    .Q(net738));
 sky130_fd_sc_hd__dlclkp_1 s869 (.CLK(clknet_4_7_0_clk),
    .GATE(net572),
    .GCLK(net739));
 sky130_fd_sc_hd__dlclkp_2 s870 (.CLK(clknet_4_7_0_clk),
    .GATE(net579),
    .GCLK(net740));
 sky130_fd_sc_hd__dlclkp_4 s871 (.CLK(clknet_4_7_0_clk),
    .GATE(net580),
    .GCLK(net741));
 sky130_fd_sc_hd__dlxbn_1 s872 (.D(net591),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net742));
 sky130_fd_sc_hd__dlxbn_1 s873 (.D(net598),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net743));
 sky130_fd_sc_hd__dlxbp_1 s874 (.D(net599),
    .GATE(clknet_4_7_0_clk),
    .Q(net745),
    .Q_N(net744));
 sky130_fd_sc_hd__dlxtn_1 s875 (.D(net601),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net746));
 sky130_fd_sc_hd__dlxtn_2 s876 (.D(net603),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net747));
 sky130_fd_sc_hd__dlxtn_1 s877 (.D(net604),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net748));
 sky130_fd_sc_hd__dlxtp_1 s878 (.D(net605),
    .GATE(clknet_4_13_0_clk),
    .Q(net749));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s879 (.D(net608),
    .SLEEP_B(clknet_4_15_0_clk),
    .Q(net750));
 sky130_fd_sc_hd__dfxbp_1 s880 (.CLK(clknet_4_15_0_clk),
    .D(net610),
    .Q(net752),
    .Q_N(net751));
 sky130_fd_sc_hd__dfxbp_1 s881 (.CLK(clknet_4_15_0_clk),
    .D(net612),
    .Q(net753));
 sky130_fd_sc_hd__dfxtp_1 s882 (.CLK(clknet_4_15_0_clk),
    .D(net616),
    .Q(net754));
 sky130_fd_sc_hd__dfxtp_1 s883 (.CLK(clknet_4_9_0_clk),
    .D(net622),
    .Q(net755));
 sky130_fd_sc_hd__dfxtp_1 s884 (.CLK(clknet_4_6_0_clk),
    .D(net623),
    .Q(net756));
 sky130_fd_sc_hd__dlclkp_1 s885 (.CLK(clknet_4_2_0_clk),
    .GATE(net636),
    .GCLK(net757));
 sky130_fd_sc_hd__dlclkp_2 s886 (.CLK(clknet_4_3_0_clk),
    .GATE(net642),
    .GCLK(net758));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net761));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_8 input5 (.A(in12),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net764));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net765));
 sky130_fd_sc_hd__buf_6 input8 (.A(in15),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in16),
    .X(net767));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(in18),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in19),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_8 input13 (.A(in2),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net772));
 sky130_fd_sc_hd__buf_2 input15 (.A(in21),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(in22),
    .X(net774));
 sky130_fd_sc_hd__buf_2 input17 (.A(in23),
    .X(net775));
 sky130_fd_sc_hd__buf_4 input18 (.A(in24),
    .X(net776));
 sky130_fd_sc_hd__buf_1 input19 (.A(in25),
    .X(net777));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(in28),
    .X(net780));
 sky130_fd_sc_hd__buf_1 input23 (.A(in29),
    .X(net781));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(in3),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net783));
 sky130_fd_sc_hd__buf_4 input26 (.A(in31),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(in33),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(in34),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(in35),
    .X(net788));
 sky130_fd_sc_hd__buf_1 input31 (.A(in36),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(in37),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(in38),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in39),
    .X(net792));
 sky130_fd_sc_hd__buf_1 input35 (.A(in4),
    .X(net793));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net794));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(in42),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net797));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net799));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net800));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in49),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(in5),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(in50),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_8 input49 (.A(in52),
    .X(net807));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(in53),
    .X(net808));
 sky130_fd_sc_hd__buf_1 input51 (.A(in54),
    .X(net809));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net810));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in57),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(in58),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net814));
 sky130_fd_sc_hd__buf_4 input57 (.A(in6),
    .X(net815));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net816));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net817));
 sky130_fd_sc_hd__buf_1 input60 (.A(in7),
    .X(net818));
 sky130_fd_sc_hd__buf_2 input61 (.A(in8),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(in9),
    .X(net820));
 sky130_fd_sc_hd__buf_2 output63 (.A(net821),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output64 (.A(net822),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net823),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(clknet_1_1__leaf_net824),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net825),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net826),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(clknet_1_1__leaf_net827),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net1015),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net829),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output72 (.A(net830),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net831),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(clknet_1_1__leaf_net832),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output75 (.A(net833),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output76 (.A(net834),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output77 (.A(net835),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output78 (.A(net836),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net837),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output80 (.A(net926),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output81 (.A(net839),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output82 (.A(net840),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output83 (.A(net841),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output84 (.A(net920),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(clknet_1_1__leaf_net843),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output86 (.A(net844),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output87 (.A(net845),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output88 (.A(net846),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output89 (.A(net847),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output90 (.A(net848),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(clknet_1_1__leaf_net849),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output92 (.A(net850),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net851),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output94 (.A(net852),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output95 (.A(net853),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output96 (.A(net929),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net855),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output98 (.A(net856),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output99 (.A(net857),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output100 (.A(net858),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(clknet_1_1__leaf_net859),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output102 (.A(net860),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output103 (.A(net861),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output104 (.A(net862),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output105 (.A(net863),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output106 (.A(net864),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output107 (.A(net865),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output108 (.A(net866),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net867),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(clknet_1_0__leaf_net868),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output111 (.A(net1030),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output112 (.A(net904),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output113 (.A(net871),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output114 (.A(net872),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output115 (.A(net873),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output116 (.A(net874),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output117 (.A(net875),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output118 (.A(net876),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output119 (.A(net877),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output120 (.A(net878),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output121 (.A(net879),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_1 max_cap122 (.A(net578),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_1 max_cap123 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_1 wire124 (.A(net539),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_1 wire125 (.A(net419),
    .X(net883));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire126 (.A(net1018),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_2 wire127 (.A(net1018),
    .X(net885));
 sky130_fd_sc_hd__buf_1 max_cap128 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__buf_1 max_cap129 (.A(net269),
    .X(net887));
 sky130_fd_sc_hd__buf_1 wire130 (.A(net225),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net890),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net362),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_2 max_cap133 (.A(net136),
    .X(net891));
 sky130_fd_sc_hd__buf_12 fanout134 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_12 fanout135 (.A(net120),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_1 max_cap136 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_1 max_cap137 (.A(net1015),
    .X(net895));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net309),
    .X(net896));
 sky130_fd_sc_hd__buf_1 max_cap139 (.A(net568),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_1 max_cap140 (.A(net424),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(net520),
    .X(net899));
 sky130_fd_sc_hd__buf_1 max_cap142 (.A(net208),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_1 max_cap143 (.A(net40),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_1 wire144 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_1 max_cap145 (.A(net299),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net870),
    .X(net904));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire147 (.A(net108),
    .X(net905));
 sky130_fd_sc_hd__buf_6 max_cap148 (.A(net108),
    .X(net906));
 sky130_fd_sc_hd__buf_1 max_cap149 (.A(net908),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_2 max_cap150 (.A(net909),
    .X(net908));
 sky130_fd_sc_hd__buf_4 max_cap151 (.A(net38),
    .X(net909));
 sky130_fd_sc_hd__buf_2 max_cap152 (.A(net263),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_1 max_cap153 (.A(net1021),
    .X(net911));
 sky130_fd_sc_hd__buf_2 max_cap154 (.A(net150),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_2 max_cap155 (.A(net36),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_2 max_cap156 (.A(net518),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net343),
    .X(net915));
 sky130_fd_sc_hd__buf_1 max_cap158 (.A(net314),
    .X(net916));
 sky130_fd_sc_hd__buf_2 wire159 (.A(net297),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__clkbuf_2 fanout161 (.A(net920),
    .X(net919));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net842),
    .X(net920));
 sky130_fd_sc_hd__buf_1 wire163 (.A(net196),
    .X(net921));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap164 (.A(net923),
    .X(net922));
 sky130_fd_sc_hd__buf_1 max_cap165 (.A(net22),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_8 fanout166 (.A(net855),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net927),
    .X(net926));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(net838),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_1 max_cap170 (.A(net78),
    .X(net928));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net854),
    .X(net929));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net729),
    .X(net930));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net695),
    .X(net931));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net696),
    .X(net932));
 sky130_fd_sc_hd__buf_6 fanout175 (.A(net767),
    .X(net933));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(net812),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net804),
    .X(net935));
 sky130_fd_sc_hd__inv_8 c556_1 (.A(clknet_1_0__leaf_net673),
    .Y(net936));
 sky130_fd_sc_hd__inv_16 c558_3 (.A(clknet_1_1__leaf_net673),
    .Y(net938));
 sky130_fd_sc_hd__inv_16 c558_4 (.A(clknet_1_0__leaf_net673),
    .Y(net939));
 sky130_fd_sc_hd__inv_16 c558_5 (.A(clknet_1_1__leaf_net673),
    .Y(net940));
 sky130_fd_sc_hd__inv_16 c558_6 (.A(clknet_1_1__leaf_net673),
    .Y(net941));
 sky130_fd_sc_hd__clkinv_1 c316_8 (.A(net675),
    .Y(net943));
 sky130_fd_sc_hd__clkinv_1 c316_9 (.A(net675),
    .Y(net944));
 sky130_fd_sc_hd__inv_12 c328_11 (.A(net675),
    .Y(net946));
 sky130_fd_sc_hd__inv_12 c328_12 (.A(net675),
    .Y(net947));
 sky130_fd_sc_hd__inv_12 c320_15 (.A(clknet_1_1__leaf_net757),
    .Y(net950));
 sky130_fd_sc_hd__inv_12 c320_16 (.A(clknet_1_0__leaf_net757),
    .Y(net951));
 sky130_fd_sc_hd__inv_12 c320_17 (.A(clknet_1_0__leaf_net757),
    .Y(net952));
 sky130_fd_sc_hd__inv_1 c449_19 (.A(clknet_1_1__leaf_net757),
    .Y(net954));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net758 (.A(net758),
    .X(clknet_0_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_0__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_1__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net431 (.A(net431),
    .X(clknet_0_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net431 (.A(clknet_0_net431),
    .X(clknet_1_0__leaf_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net431 (.A(clknet_0_net431),
    .X(clknet_1_1__leaf_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net674 (.A(net674),
    .X(clknet_0_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_1__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net465 (.A(net465),
    .X(clknet_0_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_1__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net582 (.A(net582),
    .X(clknet_0_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_0__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_1__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net611 (.A(net611),
    .X(clknet_0_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_0__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_1__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net470 (.A(net470),
    .X(clknet_0_net470));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net470 (.A(clknet_0_net470),
    .X(clknet_1_0__leaf_net470));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net470 (.A(clknet_0_net470),
    .X(clknet_1_1__leaf_net470));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net720 (.A(net720),
    .X(clknet_0_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_0__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_1__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net492 (.A(net492),
    .X(clknet_0_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_0__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_1__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net472 (.A(net472),
    .X(clknet_0_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_0__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_1__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net471 (.A(net471),
    .X(clknet_0_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_0__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_1__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net824 (.A(net824),
    .X(clknet_0_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net824 (.A(clknet_0_net824),
    .X(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net824 (.A(clknet_0_net824),
    .X(clknet_1_1__leaf_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net832 (.A(net832),
    .X(clknet_0_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net832 (.A(clknet_0_net832),
    .X(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net832 (.A(clknet_0_net832),
    .X(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net461 (.A(net461),
    .X(clknet_0_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net461 (.A(clknet_0_net461),
    .X(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net461 (.A(clknet_0_net461),
    .X(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net702 (.A(net702),
    .X(clknet_0_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_0__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_1__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net757 (.A(net757),
    .X(clknet_0_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_0__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_1__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net232 (.A(net232),
    .X(clknet_0_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net339 (.A(net339),
    .X(clknet_0_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_0__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_1__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net336 (.A(net336),
    .X(clknet_0_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_0__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_1__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net345 (.A(net345),
    .X(clknet_0_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net345 (.A(clknet_0_net345),
    .X(clknet_1_0__leaf_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net345 (.A(clknet_0_net345),
    .X(clknet_1_1__leaf_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net341 (.A(net341),
    .X(clknet_0_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_0__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_1__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net228 (.A(net228),
    .X(clknet_0_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_0__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_1__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net230 (.A(net230),
    .X(clknet_0_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net739 (.A(net739),
    .X(clknet_0_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net739 (.A(clknet_0_net739),
    .X(clknet_1_0__leaf_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net739 (.A(clknet_0_net739),
    .X(clknet_1_1__leaf_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net574 (.A(net574),
    .X(clknet_0_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_0__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_1__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net741 (.A(net741),
    .X(clknet_0_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net741 (.A(clknet_0_net741),
    .X(clknet_1_0__leaf_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net741 (.A(clknet_0_net741),
    .X(clknet_1_1__leaf_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net849 (.A(net849),
    .X(clknet_0_net849));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net849 (.A(clknet_0_net849),
    .X(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net849 (.A(clknet_0_net849),
    .X(clknet_1_1__leaf_net849));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net721 (.A(net721),
    .X(clknet_0_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_0__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_1__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net740 (.A(net740),
    .X(clknet_0_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net740 (.A(clknet_0_net740),
    .X(clknet_1_0__leaf_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net740 (.A(clknet_0_net740),
    .X(clknet_1_1__leaf_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net703 (.A(net703),
    .X(clknet_0_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net689 (.A(net689),
    .X(clknet_0_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net859 (.A(net859),
    .X(clknet_0_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net688 (.A(net688),
    .X(clknet_0_net688));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net688 (.A(clknet_0_net688),
    .X(clknet_1_0__leaf_net688));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net688 (.A(clknet_0_net688),
    .X(clknet_1_1__leaf_net688));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net687 (.A(net687),
    .X(clknet_0_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net687 (.A(clknet_0_net687),
    .X(clknet_1_0__leaf_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net687 (.A(clknet_0_net687),
    .X(clknet_1_1__leaf_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net868 (.A(net868),
    .X(clknet_0_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_1__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net827 (.A(net827),
    .X(clknet_0_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net827 (.A(clknet_0_net827),
    .X(clknet_1_0__leaf_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net827 (.A(clknet_0_net827),
    .X(clknet_1_1__leaf_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net170 (.A(net170),
    .X(clknet_0_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_0__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_1__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net673 (.A(net673),
    .X(clknet_0_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net434 (.A(net434),
    .X(clknet_0_net434));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net434 (.A(clknet_0_net434),
    .X(clknet_1_0__leaf_net434));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net434 (.A(clknet_0_net434),
    .X(clknet_1_1__leaf_net434));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net445 (.A(net445),
    .X(clknet_0_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_0__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_1__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net843 (.A(net843),
    .X(clknet_0_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net487 (.A(net487),
    .X(clknet_0_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net487 (.A(clknet_0_net487),
    .X(clknet_1_0__leaf_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net487 (.A(clknet_0_net487),
    .X(clknet_1_1__leaf_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net457 (.A(net457),
    .X(clknet_0_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_0__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_1__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net454 (.A(net454),
    .X(clknet_0_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_0__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_1__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net453 (.A(net453),
    .X(clknet_0_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net453 (.A(clknet_0_net453),
    .X(clknet_1_0__leaf_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net453 (.A(clknet_0_net453),
    .X(clknet_1_1__leaf_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net438 (.A(net438),
    .X(clknet_0_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_0__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_1__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net440 (.A(net440),
    .X(clknet_0_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_0__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_1__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net545 (.A(net545),
    .X(clknet_0_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_0__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_1__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net547 (.A(net547),
    .X(clknet_0_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net427 (.A(net427),
    .X(clknet_0_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_1__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net429 (.A(net429),
    .X(clknet_0_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_1__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net586 (.A(net586),
    .X(clknet_0_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_0__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_1__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net98),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net227),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net101),
    .X(net238));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer4 (.A(net238),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net93),
    .X(net344));
 sky130_fd_sc_hd__buf_6 rebuffer6 (.A(net112),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net426),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net426),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net108),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net956),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net223),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net958),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net959),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net960),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net961),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net961),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net119),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net964),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net213),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net213),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net967),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net79),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net969),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net893),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net971),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_1 rebuffer26 (.A(net972),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net971),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net971),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net220),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net976),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net977),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net220),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net979),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net217),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net119),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net982),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net892),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net892),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net985),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net892),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net987),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net113),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net651),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net847),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net685),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net686),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net267),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net694),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net511),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net561),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net711),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net851),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net709),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net682),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net665),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net850),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net576),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net372),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net672),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net383),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net681),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net266),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net727),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net645),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net557),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net563),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net508),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_1 wire1 (.A(net828),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(net225),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_1 max_cap3 (.A(net578),
    .X(net1017));
 sky130_fd_sc_hd__buf_1 wire4 (.A(net283),
    .X(net1018));
 sky130_fd_sc_hd__buf_1 max_cap5 (.A(net136),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_1 max_cap6 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_1 wire7 (.A(net111),
    .X(net1021));
 sky130_fd_sc_hd__buf_1 wire8 (.A(net314),
    .X(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_SCD (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SCE (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B_N (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_RESET_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_D1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_D1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_C1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_C (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A_N (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_Y (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_D (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_Y (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_D (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SET_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_SET_B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_D (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_B_N (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_C1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_Y (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_D (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_C1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_Y (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_Y (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_Y (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_SCD (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_C (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_C (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_Y (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_D1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_D (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_D (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_C_N (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_Y (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_C (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_C1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A0 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_SCD (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S0 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_X (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_C1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_C1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_RESET_B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_Y (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_C (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_C_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A_N (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Y (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_C (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B_N (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_D (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_D (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_C (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_Y (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_D1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_D (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_C (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_C (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_RESET_B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer34_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_SCD (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_RESET_B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_SCE (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_D (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_C_N (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_Y (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_RESET_B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_C_N (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_C1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net230_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_Y (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_SET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_Y (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_C_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_Y (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_SET_B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_SCD (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCE (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_D1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_C1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_D (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_S0 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_D (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_RESET_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B_N (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Y (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_C (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Y (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_D1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_C (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_Y (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_C (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_B1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_RESET_B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_C (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_C (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_SCD (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_C_N (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_SCE (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_X (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_SCE (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_D1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_Q_N (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_B_N (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_Q (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_Y (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_Q (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_C (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_C (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A_N (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_C (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_Y (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_B (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_B (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A_N (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_C_N (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_Y (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_X (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SCE (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_X (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_RESET_B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_C_N (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_X (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A3 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_Y (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_D (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_C1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_B1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_C_N (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_Y (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_Y (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_RESET_B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_Y (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_SCD (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_Q (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_Y (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_SET_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_S1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_D (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_D1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_Y (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_Q_N (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_SET_B (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold55_A (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_Q (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_SCD (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_Q_N (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B_N (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_13_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_12_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_11_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_10_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_9_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_8_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_7_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_GCLK (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_Q (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_C (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_s819_Q (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_C1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_SCD (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_s826_Q_N (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_C1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_SET_B (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_D1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_C1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_s832_Q_N (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_s832_Q (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_s834_Q (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_Q (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold53_A (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_s843_Q (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_D1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_C (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_D (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold51_A (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_Q (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_Q (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_D1 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_Q (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_D1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_Q (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_SET_B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_C1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_SET_B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_D (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A3 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_C1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_D1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_A (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_C (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_C_N (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_D_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_D1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_B1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_SCD (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A_N (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_C1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_C (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_C (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A_N (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SET_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_C (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_D1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_DE (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_B1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_C (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A3 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A_N (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_RESET_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_C1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_C (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_C (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_C (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A_N (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B_N (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A_N (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_B1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_C (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_SCE (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_C (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A_N (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_SCE (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_D1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_SCE (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_D (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_C (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B_N (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_D_N (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B_N (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_D (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_C (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_D (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_SET_B (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A_N (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_D1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_SCE (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_C (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_Y (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_C (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_D (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_Y (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_B1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_Q (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net824_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_SCE (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_B (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net832_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_RESET_B (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_Y (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_C (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_Y (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_s830_Q (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_C (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_C_N (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_D (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_Q (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net843_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_Y (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_SCE (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_SCD (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_D1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_D1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_Y (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_Y (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_s829_Q (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_D1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net849_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold52_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_Q (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_C (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_Q (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_Q (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_C_N (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_C1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_C1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_C_N (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_C (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_C (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_C_N (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_C (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_SCE (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_D1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_D (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_C (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_C_N (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCD (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_s826_Q (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_SCE (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_C (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire126_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_SCE (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_B1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer40_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer38_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer37_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_C (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap142_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_C (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_C_N (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap151_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap150_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap152_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_RESET_B (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap154_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_C1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_D (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_C1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SCD (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire159_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_C1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_D (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_C (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_S1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_C (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_C (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_C (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_D (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_C (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_C (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_X (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C_N (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_D_N (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_C (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_X (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_SCE (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_B1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SET_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_C (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_RESET_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_SCE (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_C (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_D (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_RESET_B (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_D (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_D (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SET_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_D1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_SCE (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_SCE (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_B1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_SET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_SET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_RESET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_C1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_C1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_D1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_SCE (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_D_N (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_D (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_C (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_D1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_C1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_SET_B (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_D_N (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_D1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_D (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SET_B (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_C (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_D1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_C (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_D1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_C (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B_N (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_C1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_SCD (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A_N (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_C1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_SCE (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_C_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_C (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_D (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_D (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s832_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s833_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s824_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s825_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s826_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s843_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_SLEEP_B (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s849_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s827_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s830_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s834_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s816_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s818_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s821_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s822_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s823_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_DE (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_RESET_B (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net824_X (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_SCD (.DIODE(clknet_1_1__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(clknet_1_1__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(clknet_1_1__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(clknet_1_1__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net824_X (.DIODE(clknet_1_1__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net832_A (.DIODE(clknet_0_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net832_A (.DIODE(clknet_0_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net832_X (.DIODE(clknet_0_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_SET_B (.DIODE(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCE (.DIODE(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_C (.DIODE(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net832_X (.DIODE(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A2 (.DIODE(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net832_X (.DIODE(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B_N (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_C1 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net232_X (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_SCD (.DIODE(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_SCD (.DIODE(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A1 (.DIODE(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net230_X (.DIODE(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net230_X (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net849_A (.DIODE(clknet_0_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net849_A (.DIODE(clknet_0_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net849_X (.DIODE(clknet_0_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A1 (.DIODE(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net849_X (.DIODE(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_SCE (.DIODE(clknet_1_1__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_SET_B (.DIODE(clknet_1_1__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(clknet_1_1__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_B1 (.DIODE(clknet_1_1__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(clknet_1_1__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net849_X (.DIODE(clknet_1_1__leaf_net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_C (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B1 (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net843_X (.DIODE(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net843_X (.DIODE(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C_N (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SCD (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SET_B (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_D1 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A2 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net427_X (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_C_N (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_C (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_D (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer28_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer27_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B_N (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer26_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SCE (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SET_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold53_X (.DIODE(net1000));
 sky130_fd_sc_hd__and4b_1 clone1 (.A_N(net1031),
    .B(net818),
    .C(net760),
    .D(net815),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net85),
    .X(net1024));
 sky130_fd_sc_hd__mux4_1 clone44 (.A0(net786),
    .A1(net79),
    .A2(net775),
    .A3(net780),
    .S0(net789),
    .S1(net785),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net24),
    .X(net1026));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer46 (.A(net869),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net1027),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(net1027),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net1027),
    .X(net1030));
 sky130_fd_sc_hd__buf_8 rebuffer50 (.A(net61),
    .X(net1031));
 sky130_fd_sc_hd__and3_1 clone51 (.A(net76),
    .B(net928),
    .C(net74),
    .X(net1032));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
