module netlist_4 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net750;
 wire clknet_1_0__leaf_net750;
 wire clknet_1_1__leaf_net750;
 wire clknet_0_net651;
 wire clknet_1_0__leaf_net651;
 wire clknet_1_1__leaf_net651;
 wire clknet_0_net749;
 wire clknet_1_0__leaf_net749;
 wire clknet_1_1__leaf_net749;
 wire clknet_0_net650;
 wire clknet_1_0__leaf_net650;
 wire clknet_1_1__leaf_net650;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net270;
 wire clknet_1_0__leaf_net270;
 wire clknet_1_1__leaf_net270;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net388;
 wire clknet_1_0__leaf_net388;
 wire clknet_1_1__leaf_net388;
 wire clknet_0_net500;
 wire clknet_1_0__leaf_net500;
 wire clknet_1_1__leaf_net500;
 wire clknet_0_net371;
 wire clknet_1_0__leaf_net371;
 wire clknet_1_1__leaf_net371;
 wire clknet_0_net486;
 wire clknet_1_0__leaf_net486;
 wire clknet_1_1__leaf_net486;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net581;
 wire clknet_1_0__leaf_net581;
 wire clknet_1_1__leaf_net581;
 wire clknet_0_net374;
 wire clknet_1_0__leaf_net374;
 wire clknet_1_1__leaf_net374;
 wire clknet_0_net384;
 wire clknet_1_0__leaf_net384;
 wire clknet_1_1__leaf_net384;
 wire clknet_0_net385;
 wire clknet_1_0__leaf_net385;
 wire clknet_1_1__leaf_net385;
 wire clknet_0_net377;
 wire clknet_1_0__leaf_net377;
 wire clknet_1_1__leaf_net377;
 wire clknet_0_net373;
 wire clknet_1_0__leaf_net373;
 wire clknet_1_1__leaf_net373;
 wire clknet_0_net381;
 wire clknet_1_0__leaf_net381;
 wire clknet_1_1__leaf_net381;
 wire clknet_0_net507;
 wire clknet_1_0__leaf_net507;
 wire clknet_1_1__leaf_net507;
 wire clknet_0_net513;
 wire clknet_1_0__leaf_net513;
 wire clknet_1_1__leaf_net513;
 wire clknet_0_net491;
 wire clknet_1_0__leaf_net491;
 wire clknet_1_1__leaf_net491;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net837;
 wire net840;
 wire net842;
 wire net794;
 wire net817;
 wire net836;
 wire net838;
 wire net839;
 wire net841;
 wire net843;
 wire net844;

 sky130_fd_sc_hd__o21bai_4 c100 (.A1(net45),
    .A2(net44),
    .B1_N(net35),
    .Y(net46));
 sky130_fd_sc_hd__a21boi_4 c101 (.A1(net681),
    .A2(net43),
    .B1_N(net39),
    .Y(net47));
 sky130_fd_sc_hd__and2_2 c102 (.A(net47),
    .B(net32),
    .X(net48));
 sky130_fd_sc_hd__a21bo_1 c103 (.A1(net41),
    .A2(net47),
    .B1_N(net46),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c104 (.A0(net32),
    .A1(net19),
    .A2(net7),
    .A3(net48),
    .S0(net47),
    .S1(net774),
    .X(net50));
 sky130_fd_sc_hd__nand2_1 c105 (.A(net703),
    .B(net48),
    .Y(net51));
 sky130_fd_sc_hd__nand2b_1 c106 (.A_N(net4),
    .B(net5),
    .Y(net52));
 sky130_fd_sc_hd__o21ai_1 c107 (.A1(net5),
    .A2(net48),
    .B1(net774),
    .Y(net746));
 sky130_fd_sc_hd__or2_1 c108 (.A(net51),
    .B(net11),
    .X(net53));
 sky130_fd_sc_hd__nor2b_1 c109 (.A(net746),
    .B_N(net53),
    .Y(net54));
 sky130_fd_sc_hd__or2_1 c110 (.A(net53),
    .B(net0),
    .X(net55));
 sky130_fd_sc_hd__dfrbp_1 c111 (.CLK(clknet_4_4_0_clk),
    .D(net55),
    .RESET_B(net47),
    .Q(net57),
    .Q_N(net56));
 sky130_fd_sc_hd__or2_2 c112 (.A(net708),
    .B(net53),
    .X(net58));
 sky130_fd_sc_hd__nand2_1 c113 (.A(net0),
    .B(net42),
    .Y(net59));
 sky130_fd_sc_hd__dfrbp_1 c114 (.CLK(clknet_4_4_0_clk),
    .D(net54),
    .RESET_B(net0),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__dfrtn_1 c115 (.CLK_N(clknet_4_4_0_clk),
    .D(net54),
    .RESET_B(net58),
    .Q(net62));
 sky130_fd_sc_hd__nor2_1 c116 (.A(net706),
    .B(net56),
    .Y(net63));
 sky130_fd_sc_hd__nor2_1 c117 (.A(net59),
    .B(net63),
    .Y(net64));
 sky130_fd_sc_hd__dfrtp_1 c118 (.CLK(clknet_4_4_0_clk),
    .D(net64),
    .RESET_B(net58),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_1 c119 (.CLK(clknet_4_4_0_clk),
    .D(net53),
    .RESET_B(net55),
    .Q(net66));
 sky130_fd_sc_hd__and2_2 c120 (.A(net796),
    .B(net63),
    .X(net67));
 sky130_fd_sc_hd__a21oi_1 c121 (.A1(net66),
    .A2(net60),
    .B1(net67),
    .Y(net68));
 sky130_fd_sc_hd__o31ai_1 c122 (.A1(net834),
    .A2(net68),
    .A3(net42),
    .B1(net67),
    .Y(net69));
 sky130_fd_sc_hd__a21boi_1 c123 (.A1(net57),
    .A2(net4),
    .B1_N(net67),
    .Y(net70));
 sky130_fd_sc_hd__dfbbn_1 c124 (.CLK_N(clknet_4_4_0_clk),
    .D(net69),
    .RESET_B(net11),
    .SET_B(net58),
    .Q(net731),
    .Q_N(net71));
 sky130_fd_sc_hd__dfbbn_2 c125 (.CLK_N(clknet_4_4_0_clk),
    .D(net63),
    .RESET_B(net69),
    .SET_B(net58),
    .Q(net732),
    .Q_N(net72));
 sky130_fd_sc_hd__nor2b_2 c126 (.A(net679),
    .B_N(net677),
    .Y(net73));
 sky130_fd_sc_hd__nand2b_4 c127 (.A_N(net677),
    .B(net714),
    .Y(net74));
 sky130_fd_sc_hd__or2_4 c128 (.A(net667),
    .B(net715),
    .X(net75));
 sky130_fd_sc_hd__nor2_1 c129 (.A(net73),
    .B(net677),
    .Y(net76));
 sky130_fd_sc_hd__and2_1 c130 (.A(net670),
    .B(net716),
    .X(net77));
 sky130_fd_sc_hd__or2b_2 c131 (.A(net77),
    .B_N(net700),
    .X(net78));
 sky130_fd_sc_hd__a21o_4 c132 (.A1(net675),
    .A2(net671),
    .B1(net75),
    .X(net79));
 sky130_fd_sc_hd__nor2_4 c133 (.A(net700),
    .B(net75),
    .Y(net80));
 sky130_fd_sc_hd__or2_1 c134 (.A(net79),
    .B(net668),
    .X(net81));
 sky130_fd_sc_hd__or2b_4 c135 (.A(net716),
    .B_N(net77),
    .X(net82));
 sky130_fd_sc_hd__a21oi_4 c136 (.A1(net78),
    .A2(net679),
    .B1(net82),
    .Y(net83));
 sky130_fd_sc_hd__nor2b_4 c137 (.A(net75),
    .B_N(net666),
    .Y(net84));
 sky130_fd_sc_hd__nor2_2 c138 (.A(net82),
    .B(net74),
    .Y(net85));
 sky130_fd_sc_hd__mux2_4 c139 (.A0(net80),
    .A1(net82),
    .S(net669),
    .X(net86));
 sky130_fd_sc_hd__and2_4 c140 (.A(net84),
    .B(net669),
    .X(net87));
 sky130_fd_sc_hd__mux2_4 c141 (.A0(net666),
    .A1(net85),
    .S(net87),
    .X(net88));
 sky130_fd_sc_hd__or2b_1 c142 (.A(net87),
    .B_N(net73),
    .X(net89));
 sky130_fd_sc_hd__or2b_4 c143 (.A(net89),
    .B_N(net86),
    .X(net90));
 sky130_fd_sc_hd__o41a_1 c144 (.A1(net76),
    .A2(net715),
    .A3(net90),
    .A4(net89),
    .B1(net88),
    .X(net91));
 sky130_fd_sc_hd__or2b_1 c145 (.A(net90),
    .B_N(net84),
    .X(net92));
 sky130_fd_sc_hd__nor2_4 c146 (.A(net92),
    .B(net90),
    .Y(net93));
 sky130_fd_sc_hd__nor2_1 c147 (.A(net711),
    .B(net698),
    .Y(net94));
 sky130_fd_sc_hd__nor2_2 c148 (.A(net94),
    .B(net702),
    .Y(net95));
 sky130_fd_sc_hd__or2b_1 c149 (.A(net686),
    .B_N(net671),
    .X(net96));
 sky130_fd_sc_hd__and2b_1 c150 (.A_N(net695),
    .B(net671),
    .X(net97));
 sky130_fd_sc_hd__a21o_1 c151 (.A1(net697),
    .A2(net711),
    .B1(net682),
    .X(net98));
 sky130_fd_sc_hd__nor2_2 c152 (.A(net684),
    .B(net690),
    .Y(net99));
 sky130_fd_sc_hd__nand2_2 c153 (.A(net668),
    .B(net695),
    .Y(net100));
 sky130_fd_sc_hd__nor2_1 c154 (.A(net694),
    .B(net100),
    .Y(net101));
 sky130_fd_sc_hd__nand2b_2 c155 (.A_N(net97),
    .B(net99),
    .Y(net102));
 sky130_fd_sc_hd__or2_1 c156 (.A(net102),
    .B(net101),
    .X(net103));
 sky130_fd_sc_hd__or2b_4 c157 (.A(net77),
    .B_N(net73),
    .X(net104));
 sky130_fd_sc_hd__o21a_1 c158 (.A1(net96),
    .A2(net81),
    .B1(net102),
    .X(net105));
 sky130_fd_sc_hd__or2b_1 c159 (.A(net101),
    .B_N(net102),
    .X(net106));
 sky130_fd_sc_hd__a21o_1 c160 (.A1(net84),
    .A2(net96),
    .B1(net75),
    .X(net107));
 sky130_fd_sc_hd__o31a_1 c161 (.A1(net106),
    .A2(net100),
    .A3(net97),
    .B1(net102),
    .X(net108));
 sky130_fd_sc_hd__a21o_1 c162 (.A1(net100),
    .A2(net108),
    .B1(net102),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c163 (.A0(net108),
    .A1(net102),
    .A2(net109),
    .A3(net103),
    .S0(net104),
    .S1(net106),
    .X(net110));
 sky130_fd_sc_hd__o41a_1 c164 (.A1(net97),
    .A2(net106),
    .A3(net110),
    .A4(net109),
    .B1(net94),
    .X(net111));
 sky130_fd_sc_hd__a21o_2 c165 (.A1(net105),
    .A2(net108),
    .B1(net101),
    .X(net112));
 sky130_fd_sc_hd__a21bo_1 c166 (.A1(net107),
    .A2(net110),
    .B1_N(net668),
    .X(net113));
 sky130_fd_sc_hd__and2_4 c167 (.A(net110),
    .B(net695),
    .X(net734));
 sky130_fd_sc_hd__a21oi_4 c168 (.A1(net691),
    .A2(net8),
    .B1(net773),
    .Y(net114));
 sky130_fd_sc_hd__nor2_1 c169 (.A(net114),
    .B(net717),
    .Y(net115));
 sky130_fd_sc_hd__nand2b_2 c170 (.A_N(net692),
    .B(net83),
    .Y(net116));
 sky130_fd_sc_hd__o21a_1 c171 (.A1(net2),
    .A2(net115),
    .B1(net10),
    .X(net117));
 sky130_fd_sc_hd__o21bai_4 c172 (.A1(net80),
    .A2(net114),
    .B1_N(net773),
    .Y(net118));
 sky130_fd_sc_hd__and2b_2 c173 (.A_N(net8),
    .B(net734),
    .X(net119));
 sky130_fd_sc_hd__nor2b_1 c174 (.A(net116),
    .B_N(net773),
    .Y(net120));
 sky130_fd_sc_hd__nand2_1 c175 (.A(net10),
    .B(net715),
    .Y(net121));
 sky130_fd_sc_hd__and2_2 c176 (.A(net121),
    .B(net119),
    .X(net742));
 sky130_fd_sc_hd__or2_1 c177 (.A(net115),
    .B(net773),
    .X(net122));
 sky130_fd_sc_hd__and2b_1 c178 (.A_N(net89),
    .B(net114),
    .X(net123));
 sky130_fd_sc_hd__nand2_1 c179 (.A(net123),
    .B(net103),
    .Y(net124));
 sky130_fd_sc_hd__mux2_1 c180 (.A0(net688),
    .A1(net124),
    .S(net773),
    .X(net125));
 sky130_fd_sc_hd__o21a_1 c181 (.A1(net121),
    .A2(net83),
    .B1(net119),
    .X(net126));
 sky130_fd_sc_hd__nor2_2 c182 (.A(net120),
    .B(net773),
    .Y(net127));
 sky130_fd_sc_hd__and2_1 c183 (.A(net92),
    .B(net774),
    .X(net128));
 sky130_fd_sc_hd__nor2b_2 c184 (.A(net128),
    .B_N(net123),
    .Y(net129));
 sky130_fd_sc_hd__a21o_1 c185 (.A1(net709),
    .A2(net121),
    .B1(net129),
    .X(net130));
 sky130_fd_sc_hd__nor2b_2 c186 (.A(net125),
    .B_N(net129),
    .Y(net131));
 sky130_fd_sc_hd__o21bai_4 c187 (.A1(net129),
    .A2(net131),
    .B1_N(net130),
    .Y(net132));
 sky130_fd_sc_hd__o31ai_1 c188 (.A1(net122),
    .A2(net132),
    .A3(net128),
    .B1(net119),
    .Y(net133));
 sky130_fd_sc_hd__or2b_1 c189 (.A(net690),
    .B_N(net116),
    .X(net134));
 sky130_fd_sc_hd__and2b_1 c190 (.A_N(net101),
    .B(net690),
    .X(net135));
 sky130_fd_sc_hd__and2b_1 c191 (.A_N(net130),
    .B(net698),
    .X(net136));
 sky130_fd_sc_hd__nand2_1 c192 (.A(net134),
    .B(net135),
    .Y(net137));
 sky130_fd_sc_hd__or2_4 c193 (.A(net120),
    .B(net29),
    .X(net754));
 sky130_fd_sc_hd__a21o_1 c194 (.A1(net136),
    .A2(net134),
    .B1(net83),
    .X(net138));
 sky130_fd_sc_hd__a21boi_2 c195 (.A1(net23),
    .A2(net119),
    .B1_N(net27),
    .Y(net139));
 sky130_fd_sc_hd__o41a_1 c196 (.A1(net12),
    .A2(net137),
    .A3(net134),
    .A4(net118),
    .B1(net99),
    .X(net140));
 sky130_fd_sc_hd__and2b_2 c197 (.A_N(net712),
    .B(net671),
    .X(net141));
 sky130_fd_sc_hd__nand2b_4 c198 (.A_N(net27),
    .B(net139),
    .Y(net142));
 sky130_fd_sc_hd__nor2b_1 c199 (.A(net83),
    .B_N(net140),
    .Y(net143));
 sky130_fd_sc_hd__o41a_2 c200 (.A1(net137),
    .A2(net139),
    .A3(net143),
    .A4(net141),
    .B1(net142),
    .X(net144));
 sky130_fd_sc_hd__nand2b_2 c201 (.A_N(net133),
    .B(net142),
    .Y(net145));
 sky130_fd_sc_hd__and2_1 c202 (.A(net145),
    .B(net141),
    .X(net146));
 sky130_fd_sc_hd__and2_1 c203 (.A(net143),
    .B(net138),
    .X(net147));
 sky130_fd_sc_hd__or2b_2 c204 (.A(net139),
    .B_N(net142),
    .X(net148));
 sky130_fd_sc_hd__nor2_1 c205 (.A(net17),
    .B(net137),
    .Y(net149));
 sky130_fd_sc_hd__mux2_1 c206 (.A0(net149),
    .A1(net141),
    .S(net112),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net146),
    .A1(net136),
    .A2(net149),
    .A3(net150),
    .S0(net114),
    .S1(net138),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net134),
    .A1(net140),
    .A2(net673),
    .A3(net149),
    .S0(net142),
    .S1(net151),
    .X(net152));
 sky130_fd_sc_hd__a21oi_1 c209 (.A1(net151),
    .A2(net150),
    .B1(net147),
    .Y(net153));
 sky130_fd_sc_hd__nand2_1 c210 (.A(net49),
    .B(net148),
    .Y(net154));
 sky130_fd_sc_hd__nor2b_1 c211 (.A(net33),
    .B_N(net50),
    .Y(net155));
 sky130_fd_sc_hd__nor2b_1 c212 (.A(net147),
    .B_N(net150),
    .Y(net753));
 sky130_fd_sc_hd__and2_0 c213 (.A(net116),
    .B(net144),
    .X(net156));
 sky130_fd_sc_hd__a21o_1 c214 (.A1(net39),
    .A2(net12),
    .B1(net147),
    .X(net157));
 sky130_fd_sc_hd__inv_4 c215 (.A(net639),
    .Y(net158));
 sky130_fd_sc_hd__and2b_1 c216 (.A_N(net50),
    .B(net774),
    .X(net159));
 sky130_fd_sc_hd__inv_2 c217 (.A(net638),
    .Y(net160));
 sky130_fd_sc_hd__and2b_1 c218 (.A_N(net158),
    .B(net160),
    .X(net743));
 sky130_fd_sc_hd__nand2b_1 c219 (.A_N(net160),
    .B(net158),
    .Y(net161));
 sky130_fd_sc_hd__sdfrbp_1 c220 (.CLK(clknet_4_7_0_clk),
    .D(net40),
    .RESET_B(net152),
    .SCD(net160),
    .SCE(net772),
    .Q(net163),
    .Q_N(net162));
 sky130_fd_sc_hd__a21bo_2 c221 (.A1(net15),
    .A2(net142),
    .B1_N(net157),
    .X(net739));
 sky130_fd_sc_hd__nand2b_1 c222 (.A_N(net161),
    .B(net739),
    .Y(net164));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net150),
    .A1(net141),
    .A2(net160),
    .A3(net114),
    .S0(net739),
    .S1(net157),
    .X(net165));
 sky130_fd_sc_hd__or2b_1 c224 (.A(net142),
    .B_N(net155),
    .X(net166));
 sky130_fd_sc_hd__dfbbp_1 c225 (.CLK(clknet_4_7_0_clk),
    .D(net119),
    .RESET_B(net824),
    .SET_B(net165),
    .Q(net168),
    .Q_N(net167));
 sky130_fd_sc_hd__sdfxbp_1 c226 (.CLK(clknet_4_4_0_clk),
    .D(net165),
    .SCD(net826),
    .SCE(net772),
    .Q(net170),
    .Q_N(net169));
 sky130_fd_sc_hd__mux4_2 c227 (.A0(net43),
    .A1(net772),
    .A2(net116),
    .A3(net42),
    .S0(net742),
    .S1(net159),
    .X(net171));
 sky130_fd_sc_hd__nand2_1 c228 (.A(net168),
    .B(net39),
    .Y(net172));
 sky130_fd_sc_hd__mux4_4 c229 (.A0(net171),
    .A1(net172),
    .A2(net47),
    .A3(net164),
    .S0(net33),
    .S1(net772),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net159),
    .A1(net840),
    .A2(net172),
    .A3(net772),
    .S0(net672),
    .S1(net811),
    .X(net174));
 sky130_fd_sc_hd__o21bai_1 c231 (.A1(net148),
    .A2(net46),
    .B1_N(net79),
    .Y(net175));
 sky130_fd_sc_hd__and2_1 c232 (.A(net86),
    .B(net46),
    .X(net176));
 sky130_fd_sc_hd__dfrtp_1 c233 (.CLK(clknet_4_5_0_clk),
    .D(net174),
    .RESET_B(net797),
    .Q(net177));
 sky130_fd_sc_hd__mux2_2 c234 (.A0(net176),
    .A1(net67),
    .S(net47),
    .X(net769));
 sky130_fd_sc_hd__sdfxbp_1 c235 (.CLK(clknet_4_5_0_clk),
    .D(net52),
    .SCD(net774),
    .SCE(net769),
    .Q(net179),
    .Q_N(net178));
 sky130_fd_sc_hd__dfsbp_1 c236 (.CLK(clknet_4_5_0_clk),
    .D(net140),
    .SET_B(net174),
    .Q(net181),
    .Q_N(net180));
 sky130_fd_sc_hd__or2_2 c237 (.A(net82),
    .B(net112),
    .X(net182));
 sky130_fd_sc_hd__nor2b_1 c238 (.A(net181),
    .B_N(net175),
    .Y(net183));
 sky130_fd_sc_hd__nand2b_1 c239 (.A_N(net182),
    .B(net176),
    .Y(net184));
 sky130_fd_sc_hd__and2b_1 c240 (.A_N(net177),
    .B(net732),
    .X(net185));
 sky130_fd_sc_hd__nor2_1 c241 (.A(net185),
    .B(net47),
    .Y(net718));
 sky130_fd_sc_hd__or2_1 c242 (.A(net42),
    .B(net753),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c243 (.A0(net59),
    .A1(net154),
    .A2(net718),
    .A3(net46),
    .S0(net178),
    .S1(net769),
    .X(net187));
 sky130_fd_sc_hd__o21ai_1 c244 (.A1(net185),
    .A2(net182),
    .B1(net829),
    .Y(net188));
 sky130_fd_sc_hd__sdfxtp_1 c245 (.CLK(clknet_4_4_0_clk),
    .D(net70),
    .SCD(net822),
    .SCE(net769),
    .Q(net189));
 sky130_fd_sc_hd__sdfxtp_1 c246 (.CLK(clknet_4_0_0_clk),
    .D(net814),
    .SCD(net186),
    .SCE(net183),
    .Q(net735));
 sky130_fd_sc_hd__sdfrbp_1 c247 (.CLK(clknet_4_0_0_clk),
    .D(net188),
    .RESET_B(net184),
    .SCD(net833),
    .SCE(net842),
    .Q(net191),
    .Q_N(net190));
 sky130_fd_sc_hd__o21bai_1 c248 (.A1(net175),
    .A2(net185),
    .B1_N(net70),
    .Y(net192));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net833),
    .A1(net766),
    .A2(net190),
    .A3(net742),
    .S0(net772),
    .S1(net769),
    .X(net193));
 sky130_fd_sc_hd__sdfxtp_1 c250 (.CLK(clknet_4_0_0_clk),
    .D(net769),
    .SCD(net148),
    .SCE(net819),
    .Q(net194));
 sky130_fd_sc_hd__a21boi_1 c251 (.A1(net191),
    .A2(net194),
    .B1_N(net647),
    .Y(net733));
 sky130_fd_sc_hd__nand2b_4 c252 (.A_N(net91),
    .B(net714),
    .Y(net195));
 sky130_fd_sc_hd__buf_1 c253 (.A(net73),
    .X(net196));
 sky130_fd_sc_hd__and2b_1 c254 (.A_N(net672),
    .B(net87),
    .X(net197));
 sky130_fd_sc_hd__and2_1 c255 (.A(net197),
    .B(net91),
    .X(net198));
 sky130_fd_sc_hd__inv_1 c256 (.A(net78),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 c257 (.A(net670),
    .Y(net200));
 sky130_fd_sc_hd__or2_1 c258 (.A(net200),
    .B(net88),
    .X(net201));
 sky130_fd_sc_hd__or2_1 c259 (.A(net201),
    .B(net200),
    .X(net202));
 sky130_fd_sc_hd__nor2b_1 c260 (.A(net198),
    .B_N(net201),
    .Y(net203));
 sky130_fd_sc_hd__nand2_4 c261 (.A(net202),
    .B(net200),
    .Y(net204));
 sky130_fd_sc_hd__or2_1 c262 (.A(net203),
    .B(net201),
    .X(net205));
 sky130_fd_sc_hd__nor2b_1 c263 (.A(net85),
    .B_N(net78),
    .Y(net206));
 sky130_fd_sc_hd__and2_1 c264 (.A(net205),
    .B(net206),
    .X(net207));
 sky130_fd_sc_hd__or2_2 c265 (.A(net204),
    .B(net202),
    .X(net208));
 sky130_fd_sc_hd__nor2_8 c266 (.A(net199),
    .B(net208),
    .Y(net209));
 sky130_fd_sc_hd__and2_1 c267 (.A(net202),
    .B(net204),
    .X(net210));
 sky130_fd_sc_hd__nand2b_1 c268 (.A_N(net195),
    .B(net196),
    .Y(net211));
 sky130_fd_sc_hd__nand2_1 c269 (.A(net206),
    .B(net210),
    .Y(net212));
 sky130_fd_sc_hd__o21ai_1 c270 (.A1(net210),
    .A2(net200),
    .B1(net211),
    .Y(net213));
 sky130_fd_sc_hd__or2_1 c271 (.A(net212),
    .B(net213),
    .X(net214));
 sky130_fd_sc_hd__o21bai_1 c272 (.A1(net213),
    .A2(net211),
    .B1_N(net214),
    .Y(net215));
 sky130_fd_sc_hd__or2_2 c273 (.A(net687),
    .B(net701),
    .X(net216));
 sky130_fd_sc_hd__a21boi_1 c274 (.A1(net203),
    .A2(net81),
    .B1_N(net216),
    .Y(net217));
 sky130_fd_sc_hd__or2_1 c275 (.A(net685),
    .B(net95),
    .X(net218));
 sky130_fd_sc_hd__nor2b_1 c276 (.A(net207),
    .B_N(net216),
    .Y(net219));
 sky130_fd_sc_hd__and2_4 c277 (.A(net667),
    .B(net200),
    .X(net220));
 sky130_fd_sc_hd__or2b_1 c278 (.A(net693),
    .B_N(net98),
    .X(net221));
 sky130_fd_sc_hd__nor2_1 c279 (.A(net221),
    .B(net220),
    .Y(net222));
 sky130_fd_sc_hd__and2b_1 c280 (.A_N(net214),
    .B(net113),
    .X(net223));
 sky130_fd_sc_hd__or2b_4 c281 (.A(net220),
    .B_N(net88),
    .X(net224));
 sky130_fd_sc_hd__and2_1 c282 (.A(net219),
    .B(net223),
    .X(net225));
 sky130_fd_sc_hd__nor2b_1 c283 (.A(net222),
    .B_N(net109),
    .Y(net226));
 sky130_fd_sc_hd__nor2_1 c284 (.A(net81),
    .B(net222),
    .Y(net227));
 sky130_fd_sc_hd__or2_1 c285 (.A(net217),
    .B(net81),
    .X(net228));
 sky130_fd_sc_hd__o31a_1 c286 (.A1(net219),
    .A2(net207),
    .A3(net227),
    .B1(net224),
    .X(net229));
 sky130_fd_sc_hd__nand2_1 c287 (.A(net229),
    .B(net224),
    .Y(net230));
 sky130_fd_sc_hd__o31ai_1 c288 (.A1(net227),
    .A2(net214),
    .A3(net230),
    .B1(net224),
    .Y(net231));
 sky130_fd_sc_hd__and2_1 c289 (.A(net227),
    .B(net770),
    .X(net232));
 sky130_fd_sc_hd__o21bai_1 c290 (.A1(net231),
    .A2(net230),
    .B1_N(net770),
    .Y(net233));
 sky130_fd_sc_hd__sdfbbn_1 c291 (.CLK_N(clknet_4_9_0_clk),
    .D(net226),
    .RESET_B(net734),
    .SCD(net233),
    .SCE(net770),
    .SET_B(net98),
    .Q(net235),
    .Q_N(net234));
 sky130_fd_sc_hd__and2_4 c292 (.A(net224),
    .B(net197),
    .X(net236));
 sky130_fd_sc_hd__dfsbp_1 c293 (.CLK(clknet_4_9_0_clk),
    .D(net233),
    .SET_B(net236),
    .Q(net238),
    .Q_N(net237));
 sky130_fd_sc_hd__nor2_1 c294 (.A(net717),
    .B(net770),
    .Y(net239));
 sky130_fd_sc_hd__o21ba_1 c295 (.A1(net126),
    .A2(net223),
    .B1_N(net88),
    .X(net240));
 sky130_fd_sc_hd__and2b_1 c296 (.A_N(net239),
    .B(net131),
    .X(net241));
 sky130_fd_sc_hd__nand2b_1 c297 (.A_N(net240),
    .B(net770),
    .Y(net242));
 sky130_fd_sc_hd__nor2_1 c298 (.A(net128),
    .B(net126),
    .Y(net243));
 sky130_fd_sc_hd__or2b_1 c299 (.A(net200),
    .B_N(net242),
    .X(net244));
 sky130_fd_sc_hd__nor2_1 c300 (.A(net241),
    .B(net118),
    .Y(net245));
 sky130_fd_sc_hd__and2_0 c301 (.A(net222),
    .B(net200),
    .X(net246));
 sky130_fd_sc_hd__or2_2 c302 (.A(net131),
    .B(net242),
    .X(net247));
 sky130_fd_sc_hd__nand2_1 c303 (.A(net123),
    .B(net223),
    .Y(net248));
 sky130_fd_sc_hd__and2_1 c304 (.A(net230),
    .B(net242),
    .X(net249));
 sky130_fd_sc_hd__and2_1 c305 (.A(net223),
    .B(net200),
    .X(net250));
 sky130_fd_sc_hd__a21oi_1 c306 (.A1(net246),
    .A2(net249),
    .B1(net126),
    .Y(net251));
 sky130_fd_sc_hd__and2_4 c307 (.A(net247),
    .B(net100),
    .X(net252));
 sky130_fd_sc_hd__nand2_4 c308 (.A(net250),
    .B(net240),
    .Y(net758));
 sky130_fd_sc_hd__mux4_4 c309 (.A0(net243),
    .A1(net200),
    .A2(net252),
    .A3(net245),
    .S0(net682),
    .S1(net223),
    .X(net253));
 sky130_fd_sc_hd__nand2_1 c310 (.A(net244),
    .B(net247),
    .Y(net254));
 sky130_fd_sc_hd__nand2_1 c311 (.A(net129),
    .B(net758),
    .Y(net255));
 sky130_fd_sc_hd__dfstp_1 c312 (.CLK(clknet_4_9_0_clk),
    .D(net251),
    .SET_B(net222),
    .Q(net256));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net256),
    .A1(net249),
    .A2(net251),
    .A3(net240),
    .S0(net252),
    .S1(net648),
    .X(net257));
 sky130_fd_sc_hd__dfstp_1 c314 (.CLK(clknet_4_9_0_clk),
    .D(net251),
    .SET_B(net795),
    .Q(net258));
 sky130_fd_sc_hd__nand2b_2 c315 (.A_N(net248),
    .B(net138),
    .Y(net259));
 sky130_fd_sc_hd__o31a_1 c316 (.A1(net704),
    .A2(net114),
    .A3(net258),
    .B1(net774),
    .X(net260));
 sky130_fd_sc_hd__nor2_4 c317 (.A(net220),
    .B(net648),
    .Y(net740));
 sky130_fd_sc_hd__mux2_1 c318 (.A0(net701),
    .A1(net114),
    .S(net682),
    .X(net261));
 sky130_fd_sc_hd__nand2b_1 c319 (.A_N(net260),
    .B(net831),
    .Y(net262));
 sky130_fd_sc_hd__dfbbn_1 c320 (.CLK_N(clknet_4_6_0_clk),
    .D(net153),
    .RESET_B(net95),
    .SET_B(net770),
    .Q(net264),
    .Q_N(net263));
 sky130_fd_sc_hd__o21ai_2 c321 (.A1(net138),
    .A2(net770),
    .B1(net263),
    .Y(net265));
 sky130_fd_sc_hd__a21bo_1 c322 (.A1(net677),
    .A2(net263),
    .B1_N(net837),
    .X(net266));
 sky130_fd_sc_hd__o21ai_4 c323 (.A1(net266),
    .A2(net24),
    .B1(net247),
    .Y(net267));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net74),
    .A1(net267),
    .A2(net259),
    .A3(net138),
    .S0(net698),
    .S1(net648),
    .X(net268));
 sky130_fd_sc_hd__mux4_4 c325 (.A0(net1),
    .A1(net264),
    .A2(net758),
    .A3(net204),
    .S0(net740),
    .S1(clknet_1_1__leaf_net650),
    .X(net269));
 sky130_fd_sc_hd__and2b_2 c326 (.A_N(clknet_1_0__leaf_net269),
    .B(net839),
    .X(net270));
 sky130_fd_sc_hd__and2_1 c327 (.A(net261),
    .B(net740),
    .X(net271));
 sky130_fd_sc_hd__nand2_4 c328 (.A(net271),
    .B(net259),
    .Y(net765));
 sky130_fd_sc_hd__dfbbn_1 c329 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net270),
    .RESET_B(net247),
    .SET_B(net765),
    .Q(net272));
 sky130_fd_sc_hd__o21ba_2 c330 (.A1(net264),
    .A2(clknet_1_1__leaf_net269),
    .B1_N(net265),
    .X(net273));
 sky130_fd_sc_hd__o21ba_1 c331 (.A1(net262),
    .A2(net264),
    .B1_N(net765),
    .X(net274));
 sky130_fd_sc_hd__dfbbp_1 c332 (.CLK(clknet_4_12_0_clk),
    .D(net715),
    .RESET_B(clknet_1_0__leaf_net270),
    .SET_B(net267),
    .Q(net276),
    .Q_N(net275));
 sky130_fd_sc_hd__dfstp_4 c333 (.CLK(clknet_4_2_0_clk),
    .D(net274),
    .SET_B(clknet_1_0__leaf_net650),
    .Q(net768));
 sky130_fd_sc_hd__a21bo_1 c334 (.A1(net272),
    .A2(net768),
    .B1_N(net765),
    .X(net277));
 sky130_fd_sc_hd__mux4_2 c335 (.A0(net274),
    .A1(net21),
    .A2(net204),
    .A3(net765),
    .S0(net144),
    .S1(clknet_1_1__leaf_net270),
    .X(net278));
 sky130_fd_sc_hd__dlrbn_1 c336 (.D(net164),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net112),
    .Q(net280),
    .Q_N(net279));
 sky130_fd_sc_hd__nand2b_1 c337 (.A_N(net163),
    .B(net204),
    .Y(net281));
 sky130_fd_sc_hd__and2b_1 c338 (.A_N(net172),
    .B(net279),
    .X(net282));
 sky130_fd_sc_hd__and2_1 c339 (.A(net170),
    .B(net104),
    .X(net283));
 sky130_fd_sc_hd__or2b_1 c340 (.A(net31),
    .B_N(net144),
    .X(net284));
 sky130_fd_sc_hd__and2_0 c341 (.A(net144),
    .B(net118),
    .X(net285));
 sky130_fd_sc_hd__sdfxbp_1 c342 (.CLK(clknet_4_7_0_clk),
    .D(net284),
    .SCD(net265),
    .SCE(net164),
    .Q(net286));
 sky130_fd_sc_hd__nand2_1 c343 (.A(net285),
    .B(net74),
    .Y(net287));
 sky130_fd_sc_hd__nor2b_1 c344 (.A(net770),
    .B_N(net739),
    .Y(net288));
 sky130_fd_sc_hd__nor2_1 c345 (.A(net156),
    .B(net287),
    .Y(net289));
 sky130_fd_sc_hd__and2b_1 c346 (.A_N(net289),
    .B(net281),
    .X(net290));
 sky130_fd_sc_hd__and2b_1 c347 (.A_N(net157),
    .B(net209),
    .X(net291));
 sky130_fd_sc_hd__and2_0 c348 (.A(net45),
    .B(net770),
    .X(net292));
 sky130_fd_sc_hd__o31ai_1 c349 (.A1(net828),
    .A2(net48),
    .A3(net38),
    .B1(net770),
    .Y(net293));
 sky130_fd_sc_hd__sdfbbn_1 c350 (.CLK_N(clknet_4_2_0_clk),
    .D(net293),
    .RESET_B(net288),
    .SCD(net156),
    .SCE(net768),
    .SET_B(net740),
    .Q(net294));
 sky130_fd_sc_hd__dlrbn_1 c351 (.D(net288),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net45),
    .Q(net296),
    .Q_N(net295));
 sky130_fd_sc_hd__nor2b_1 c352 (.A(net294),
    .B_N(net296),
    .Y(net297));
 sky130_fd_sc_hd__o41a_4 c353 (.A1(net291),
    .A2(net161),
    .A3(net836),
    .A4(net827),
    .B1(net46),
    .X(net298));
 sky130_fd_sc_hd__sdfxbp_1 c354 (.CLK(clknet_4_1_0_clk),
    .D(net282),
    .SCD(net298),
    .SCE(net161),
    .Q(net300),
    .Q_N(net299));
 sky130_fd_sc_hd__sdfxtp_1 c355 (.CLK(clknet_4_1_0_clk),
    .D(net812),
    .SCD(net297),
    .SCE(net298),
    .Q(net301));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net301),
    .A1(net225),
    .A2(net295),
    .A3(net291),
    .S0(net284),
    .S1(net768),
    .X(net302));
 sky130_fd_sc_hd__a21boi_0 c357 (.A1(net283),
    .A2(net104),
    .B1_N(net758),
    .Y(net303));
 sky130_fd_sc_hd__a21boi_1 c358 (.A1(net259),
    .A2(net296),
    .B1_N(net810),
    .Y(net304));
 sky130_fd_sc_hd__sdfxtp_1 c359 (.CLK(clknet_4_4_0_clk),
    .D(net48),
    .SCD(net298),
    .SCE(net60),
    .Q(net305));
 sky130_fd_sc_hd__dlrbp_1 c360 (.D(net183),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net772),
    .Q(net307),
    .Q_N(net306));
 sky130_fd_sc_hd__dlrbp_1 c361 (.D(net184),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net177),
    .Q(net308));
 sky130_fd_sc_hd__dlrtn_1 c362 (.D(net192),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net798),
    .Q(net309));
 sky130_fd_sc_hd__a21oi_1 c363 (.A1(net68),
    .A2(net303),
    .B1(net827),
    .Y(net310));
 sky130_fd_sc_hd__nor2_1 c364 (.A(net305),
    .B(net71),
    .Y(net311));
 sky130_fd_sc_hd__a21bo_1 c365 (.A1(net308),
    .A2(net61),
    .B1_N(net306),
    .X(net312));
 sky130_fd_sc_hd__sdfxtp_1 c366 (.CLK(clknet_4_0_0_clk),
    .D(net154),
    .SCD(net769),
    .SCE(net774),
    .Q(net757));
 sky130_fd_sc_hd__a21boi_1 c367 (.A1(net671),
    .A2(net194),
    .B1_N(net774),
    .Y(net313));
 sky130_fd_sc_hd__a21boi_1 c368 (.A1(net713),
    .A2(net311),
    .B1_N(net754),
    .Y(net314));
 sky130_fd_sc_hd__dfbbn_1 c369 (.CLK_N(clknet_4_5_0_clk),
    .D(net67),
    .RESET_B(net310),
    .SET_B(net61),
    .Q(net315));
 sky130_fd_sc_hd__o21bai_1 c370 (.A1(net61),
    .A2(net798),
    .B1_N(net810),
    .Y(net316));
 sky130_fd_sc_hd__dlrtn_1 c371 (.D(net58),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net316),
    .Q(net317));
 sky130_fd_sc_hd__or2b_1 c372 (.A(net292),
    .B_N(net315),
    .X(net756));
 sky130_fd_sc_hd__o21bai_2 c373 (.A1(net112),
    .A2(net317),
    .B1_N(net758),
    .Y(net318));
 sky130_fd_sc_hd__o31a_1 c374 (.A1(net314),
    .A2(net318),
    .A3(net732),
    .B1(net209),
    .X(net319));
 sky130_fd_sc_hd__sdfrtn_1 c375 (.CLK_N(clknet_4_5_0_clk),
    .D(net319),
    .RESET_B(net312),
    .SCD(net772),
    .SCE(net757),
    .Q(net320));
 sky130_fd_sc_hd__dfbbn_1 c376 (.CLK_N(clknet_4_5_0_clk),
    .D(net313),
    .RESET_B(net800),
    .SET_B(net319),
    .Q(net322),
    .Q_N(net321));
 sky130_fd_sc_hd__o31ai_1 c377 (.A1(net317),
    .A2(net318),
    .A3(net718),
    .B1(net316),
    .Y(net747));
 sky130_fd_sc_hd__or2_1 c378 (.A(net215),
    .B(net198),
    .X(net323));
 sky130_fd_sc_hd__and2_1 c379 (.A(net675),
    .B(net211),
    .X(net324));
 sky130_fd_sc_hd__nor2_1 c380 (.A(net211),
    .B(net215),
    .Y(net325));
 sky130_fd_sc_hd__nand2b_2 c381 (.A_N(net90),
    .B(net93),
    .Y(net326));
 sky130_fd_sc_hd__and2_1 c382 (.A(net326),
    .B(net79),
    .X(net327));
 sky130_fd_sc_hd__and2_2 c383 (.A(net323),
    .B(net326),
    .X(net328));
 sky130_fd_sc_hd__and2_1 c384 (.A(net327),
    .B(net326),
    .X(net329));
 sky130_fd_sc_hd__and2_1 c385 (.A(net323),
    .B(net673),
    .X(net330));
 sky130_fd_sc_hd__or2b_1 c386 (.A(net329),
    .B_N(net330),
    .X(net331));
 sky130_fd_sc_hd__or2_1 c387 (.A(net330),
    .B(net328),
    .X(net332));
 sky130_fd_sc_hd__inv_1 c388 (.A(net196),
    .Y(net333));
 sky130_fd_sc_hd__nor2b_1 c389 (.A(net333),
    .B_N(net332),
    .Y(net334));
 sky130_fd_sc_hd__mux2_1 c390 (.A0(net327),
    .A1(net324),
    .S(net211),
    .X(net335));
 sky130_fd_sc_hd__and2_1 c391 (.A(net331),
    .B(net196),
    .X(net336));
 sky130_fd_sc_hd__and2b_1 c392 (.A_N(net325),
    .B(net333),
    .X(net337));
 sky130_fd_sc_hd__and2_1 c393 (.A(net331),
    .B(net332),
    .X(net338));
 sky130_fd_sc_hd__nor2_4 c394 (.A(net335),
    .B(net328),
    .Y(net339));
 sky130_fd_sc_hd__sdfbbp_1 c395 (.CLK(clknet_4_8_0_clk),
    .D(net330),
    .RESET_B(net336),
    .SCD(net338),
    .SCE(net339),
    .SET_B(net333),
    .Q(net341),
    .Q_N(net340));
 sky130_fd_sc_hd__dlrtn_1 c396 (.D(net334),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net801),
    .Q(net342));
 sky130_fd_sc_hd__dlrtp_2 c397 (.D(net338),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net330),
    .Q(net343));
 sky130_fd_sc_hd__or2_4 c398 (.A(net341),
    .B(net328),
    .X(net751));
 sky130_fd_sc_hd__and2b_2 c399 (.A_N(net235),
    .B(net104),
    .X(net344));
 sky130_fd_sc_hd__and2_1 c400 (.A(net208),
    .B(net751),
    .X(net345));
 sky130_fd_sc_hd__nand2_4 c401 (.A(net236),
    .B(net237),
    .Y(net346));
 sky130_fd_sc_hd__and2b_1 c402 (.A_N(net342),
    .B(net226),
    .X(net347));
 sky130_fd_sc_hd__or2_4 c403 (.A(net218),
    .B(net346),
    .X(net752));
 sky130_fd_sc_hd__dlrtp_1 c404 (.D(net344),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net345),
    .Q(net348));
 sky130_fd_sc_hd__dlrtp_1 c405 (.D(net224),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net345),
    .Q(net349));
 sky130_fd_sc_hd__dfbbp_1 c406 (.CLK(clknet_4_8_0_clk),
    .D(net345),
    .RESET_B(net234),
    .SET_B(net804),
    .Q(net351),
    .Q_N(net350));
 sky130_fd_sc_hd__and2b_1 c407 (.A_N(net348),
    .B(net195),
    .X(net352));
 sky130_fd_sc_hd__or2_4 c408 (.A(net109),
    .B(net752),
    .X(net353));
 sky130_fd_sc_hd__a21bo_1 c409 (.A1(net75),
    .A2(net353),
    .B1_N(net347),
    .X(net354));
 sky130_fd_sc_hd__and2_1 c410 (.A(net98),
    .B(net350),
    .X(net355));
 sky130_fd_sc_hd__and2_2 c411 (.A(net353),
    .B(net347),
    .X(net356));
 sky130_fd_sc_hd__nand2b_1 c412 (.A_N(net346),
    .B(net344),
    .Y(net357));
 sky130_fd_sc_hd__mux2_4 c413 (.A0(net351),
    .A1(net226),
    .S(net216),
    .X(net358));
 sky130_fd_sc_hd__o41a_4 c414 (.A1(net358),
    .A2(net351),
    .A3(net352),
    .A4(net353),
    .B1(net780),
    .X(net359));
 sky130_fd_sc_hd__edfxbp_1 c415 (.CLK(clknet_4_8_0_clk),
    .D(net336),
    .DE(net356),
    .Q(net361),
    .Q_N(net360));
 sky130_fd_sc_hd__nor2_4 c416 (.A(net228),
    .B(net359),
    .Y(net362));
 sky130_fd_sc_hd__o21bai_4 c417 (.A1(net356),
    .A2(net789),
    .B1_N(net357),
    .Y(net363));
 sky130_fd_sc_hd__sdfbbn_1 c418 (.CLK_N(clknet_4_8_0_clk),
    .D(net349),
    .RESET_B(net345),
    .SCD(net815),
    .SCE(net358),
    .SET_B(net752),
    .Q(net364));
 sky130_fd_sc_hd__o21ba_1 c419 (.A1(net357),
    .A2(net364),
    .B1_N(net358),
    .X(net365));
 sky130_fd_sc_hd__a21boi_1 c420 (.A1(net790),
    .A2(net359),
    .B1_N(net242),
    .Y(net366));
 sky130_fd_sc_hd__a21o_2 c421 (.A1(net698),
    .A2(net220),
    .B1(net784),
    .X(net367));
 sky130_fd_sc_hd__a21bo_1 c422 (.A1(net357),
    .A2(net355),
    .B1_N(net698),
    .X(net368));
 sky130_fd_sc_hd__or2_1 c423 (.A(net676),
    .B(net220),
    .X(net369));
 sky130_fd_sc_hd__edfxtp_1 c424 (.CLK(clknet_4_9_0_clk),
    .D(net254),
    .DE(net220),
    .Q(net370));
 sky130_fd_sc_hd__sdlclkp_1 c425 (.CLK(clknet_4_6_0_clk),
    .GATE(net245),
    .SCE(net103),
    .GCLK(net371));
 sky130_fd_sc_hd__nand2_1 c426 (.A(net240),
    .B(net99),
    .Y(net372));
 sky130_fd_sc_hd__or2b_4 c427 (.A(net362),
    .B_N(clknet_1_0__leaf_net371),
    .X(net373));
 sky130_fd_sc_hd__a21oi_2 c428 (.A1(clknet_1_1__leaf_net373),
    .A2(clknet_1_0__leaf_net371),
    .B1(net367),
    .Y(net374));
 sky130_fd_sc_hd__or2_1 c429 (.A(net249),
    .B(net368),
    .X(net375));
 sky130_fd_sc_hd__o21ba_1 c430 (.A1(net365),
    .A2(net117),
    .B1_N(net362),
    .X(net376));
 sky130_fd_sc_hd__or2_4 c431 (.A(clknet_1_1__leaf_net374),
    .B(net361),
    .X(net377));
 sky130_fd_sc_hd__and2b_1 c432 (.A_N(net366),
    .B(net359),
    .X(net378));
 sky130_fd_sc_hd__sdfxbp_1 c433 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net374),
    .SCD(net348),
    .SCE(net378),
    .Q(net380),
    .Q_N(net379));
 sky130_fd_sc_hd__o21ba_4 c434 (.A1(net370),
    .A2(net195),
    .B1_N(net369),
    .X(net744));
 sky130_fd_sc_hd__o21ai_4 c435 (.A1(net356),
    .A2(clknet_1_0__leaf_net373),
    .B1(net370),
    .Y(net381));
 sky130_fd_sc_hd__sdfbbn_1 c436 (.CLK_N(clknet_4_9_0_clk),
    .D(net786),
    .RESET_B(net378),
    .SCD(net375),
    .SCE(net791),
    .SET_B(clknet_1_0__leaf_net381),
    .Q(net383),
    .Q_N(net382));
 sky130_fd_sc_hd__o41a_2 c437 (.A1(net368),
    .A2(net702),
    .A3(net383),
    .A4(clknet_1_0__leaf_net374),
    .B1(net367),
    .X(net384));
 sky130_fd_sc_hd__a21boi_2 c438 (.A1(net380),
    .A2(clknet_1_0__leaf_net384),
    .B1_N(net383),
    .Y(net385));
 sky130_fd_sc_hd__sdfrtp_1 c439 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net385),
    .RESET_B(clknet_1_0__leaf_net371),
    .SCD(net379),
    .SCE(clknet_1_0__leaf_net384),
    .Q(net386));
 sky130_fd_sc_hd__sdfxbp_1 c440 (.CLK(clknet_4_12_0_clk),
    .D(net255),
    .SCD(clknet_1_0__leaf_net385),
    .SCE(clknet_1_0__leaf_net381),
    .Q(net387));
 sky130_fd_sc_hd__sdlclkp_2 c441 (.CLK(clknet_4_7_0_clk),
    .GATE(net837),
    .SCE(net277),
    .GCLK(net388));
 sky130_fd_sc_hd__sdlclkp_4 c442 (.CLK(clknet_4_12_0_clk),
    .GATE(net265),
    .SCE(net375),
    .GCLK(net389));
 sky130_fd_sc_hd__nand2_1 c443 (.A(net673),
    .B(clknet_1_1__leaf_net381),
    .Y(net390));
 sky130_fd_sc_hd__or2b_2 c444 (.A(net29),
    .B_N(net768),
    .X(net391));
 sky130_fd_sc_hd__nand2b_1 c445 (.A_N(net386),
    .B(net24),
    .Y(net392));
 sky130_fd_sc_hd__nand2b_1 c446 (.A_N(net387),
    .B(net391),
    .Y(net393));
 sky130_fd_sc_hd__nand2_1 c447 (.A(net393),
    .B(net363),
    .Y(net394));
 sky130_fd_sc_hd__sdfbbp_1 c448 (.CLK(clknet_4_7_0_clk),
    .D(net394),
    .RESET_B(net754),
    .SCD(net220),
    .SCE(net252),
    .SET_B(net391),
    .Q(net396),
    .Q_N(net395));
 sky130_fd_sc_hd__o21ai_0 c449 (.A1(net276),
    .A2(net339),
    .B1(net145),
    .Y(net397));
 sky130_fd_sc_hd__nor2_2 c450 (.A(net391),
    .B(clknet_1_0__leaf_net651),
    .Y(net398));
 sky130_fd_sc_hd__sdfrtp_4 c451 (.CLK(clknet_4_2_0_clk),
    .D(net397),
    .RESET_B(net274),
    .SCD(net275),
    .SCE(net391),
    .Q(net729));
 sky130_fd_sc_hd__sdfrtp_1 c452 (.CLK(clknet_4_2_0_clk),
    .D(net376),
    .RESET_B(net252),
    .SCD(net394),
    .SCE(net28),
    .Q(net399));
 sky130_fd_sc_hd__or2_1 c453 (.A(net220),
    .B(net396),
    .X(net759));
 sky130_fd_sc_hd__o21ba_2 c454 (.A1(net95),
    .A2(clknet_1_1__leaf_net388),
    .B1_N(net729),
    .X(net400));
 sky130_fd_sc_hd__nand2b_1 c455 (.A_N(net391),
    .B(clknet_1_1__leaf_net651),
    .Y(net401));
 sky130_fd_sc_hd__nor2_1 c456 (.A(net400),
    .B(net95),
    .Y(net738));
 sky130_fd_sc_hd__dfrbp_1 c457 (.CLK(clknet_4_7_0_clk),
    .D(net273),
    .RESET_B(net729),
    .Q(net402));
 sky130_fd_sc_hd__nor2_1 c458 (.A(net399),
    .B(net401),
    .Y(net403));
 sky130_fd_sc_hd__o21ba_2 c459 (.A1(net403),
    .A2(net382),
    .B1_N(net395),
    .X(net404));
 sky130_fd_sc_hd__mux4_2 c460 (.A0(net398),
    .A1(net265),
    .A2(net386),
    .A3(net220),
    .S0(net794),
    .S1(clknet_1_0__leaf_net388),
    .X(net749));
 sky130_fd_sc_hd__nor2_2 c461 (.A(net404),
    .B(clknet_1_0__leaf_net749),
    .Y(net405));
 sky130_fd_sc_hd__and2b_4 c462 (.A_N(net99),
    .B(net754),
    .X(net406));
 sky130_fd_sc_hd__or2b_1 c463 (.A(net38),
    .B_N(net775),
    .X(net407));
 sky130_fd_sc_hd__o21bai_4 c464 (.A1(net744),
    .A2(net754),
    .B1_N(net645),
    .Y(net408));
 sky130_fd_sc_hd__clkbuf_1 c465 (.A(net665),
    .X(net409));
 sky130_fd_sc_hd__nor2_1 c466 (.A(net369),
    .B(net406),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 c467 (.A(net665),
    .Y(net411));
 sky130_fd_sc_hd__sdfbbn_1 c468 (.CLK_N(clknet_4_2_0_clk),
    .D(net302),
    .RESET_B(net369),
    .SCD(clknet_1_0__leaf_net749),
    .SCE(net395),
    .SET_B(net408),
    .Q(net412));
 sky130_fd_sc_hd__o21ba_1 c469 (.A1(net104),
    .A2(net406),
    .B1_N(net339),
    .X(net760));
 sky130_fd_sc_hd__o21ai_1 c470 (.A1(net396),
    .A2(net765),
    .B1(net209),
    .Y(net413));
 sky130_fd_sc_hd__sdfxtp_1 c471 (.CLK(clknet_4_2_0_clk),
    .D(net408),
    .SCD(net290),
    .SCE(net298),
    .Q(net414));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net411),
    .A1(net408),
    .A2(net413),
    .A3(net765),
    .S0(net406),
    .S1(net739),
    .X(net415));
 sky130_fd_sc_hd__and2_1 c473 (.A(net412),
    .B(net406),
    .X(net416));
 sky130_fd_sc_hd__sdfxtp_1 c474 (.CLK(clknet_4_3_0_clk),
    .D(net413),
    .SCD(net820),
    .SCE(clknet_1_0__leaf_net388),
    .Q(net417));
 sky130_fd_sc_hd__o21ai_1 c475 (.A1(net414),
    .A2(net408),
    .B1(net396),
    .Y(net418));
 sky130_fd_sc_hd__a21oi_1 c476 (.A1(net416),
    .A2(net408),
    .B1(net410),
    .Y(net419));
 sky130_fd_sc_hd__o21ai_4 c477 (.A1(net406),
    .A2(net417),
    .B1(net652),
    .Y(net750));
 sky130_fd_sc_hd__o41a_1 c478 (.A1(net409),
    .A2(net406),
    .A3(net417),
    .A4(net772),
    .B1(net739),
    .X(net420));
 sky130_fd_sc_hd__or2b_2 c479 (.A(net402),
    .B_N(net419),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net390),
    .A1(net418),
    .A2(net410),
    .A3(net421),
    .S0(net413),
    .S1(net414),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net417),
    .A1(net421),
    .A2(net408),
    .A3(net298),
    .S0(net406),
    .S1(net653),
    .X(net423));
 sky130_fd_sc_hd__o31ai_4 c482 (.A1(net410),
    .A2(net421),
    .A3(net339),
    .B1(net654),
    .Y(net424));
 sky130_fd_sc_hd__o31ai_1 c494 (.A1(net296),
    .A2(net307),
    .A3(net758),
    .B1(net318),
    .Y(net425));
 sky130_fd_sc_hd__sdfsbp_1 c495 (.CLK(clknet_4_1_0_clk),
    .D(net298),
    .SCD(net209),
    .SCE(net104),
    .SET_B(net72),
    .Q(net745));
 sky130_fd_sc_hd__o41a_2 c496 (.A1(net186),
    .A2(net311),
    .A3(net79),
    .A4(net807),
    .B1(net304),
    .X(net764));
 sky130_fd_sc_hd__sdfbbn_1 c497 (.CLK_N(clknet_4_0_0_clk),
    .D(net813),
    .RESET_B(net304),
    .SCD(net267),
    .SCE(net765),
    .SET_B(net298),
    .Q(net426));
 sky130_fd_sc_hd__o31ai_1 c498 (.A1(net300),
    .A2(net756),
    .A3(net307),
    .B1(net72),
    .Y(net724));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net118),
    .A1(net318),
    .A2(net46),
    .A3(net744),
    .S0(net756),
    .S1(net772),
    .X(net723));
 sky130_fd_sc_hd__sdfbbp_1 c500 (.CLK(clknet_4_0_0_clk),
    .D(net267),
    .RESET_B(net807),
    .SCD(net321),
    .SCE(net817),
    .SET_B(net802),
    .Q(net761));
 sky130_fd_sc_hd__sdfbbn_1 c501 (.CLK_N(clknet_4_1_0_clk),
    .D(net818),
    .RESET_B(net808),
    .SCD(net757),
    .SCE(net764),
    .SET_B(net420),
    .Q(net762));
 sky130_fd_sc_hd__sdfsbp_1 c502 (.CLK(clknet_4_1_0_clk),
    .D(net425),
    .SCD(net186),
    .SCE(net72),
    .SET_B(net764),
    .Q(net755));
 sky130_fd_sc_hd__sdfbbn_1 c503 (.CLK_N(clknet_4_1_0_clk),
    .D(net46),
    .RESET_B(net420),
    .SCD(net754),
    .SCE(net299),
    .SET_B(net776),
    .Q(net730));
 sky130_fd_sc_hd__clkbuf_1 c504 (.A(net689),
    .X(net427));
 sky130_fd_sc_hd__nor2b_1 c505 (.A(net87),
    .B_N(net751),
    .Y(net428));
 sky130_fd_sc_hd__clkbuf_2 c506 (.A(net212),
    .X(net429));
 sky130_fd_sc_hd__nand2b_1 c507 (.A_N(net717),
    .B(net87),
    .Y(net430));
 sky130_fd_sc_hd__or2b_2 c508 (.A(net85),
    .B_N(net93),
    .X(net431));
 sky130_fd_sc_hd__and2b_1 c509 (.A_N(net430),
    .B(net76),
    .X(net432));
 sky130_fd_sc_hd__nor2b_4 c510 (.A(net328),
    .B_N(net327),
    .Y(net433));
 sky130_fd_sc_hd__and2_1 c511 (.A(net427),
    .B(net433),
    .X(net434));
 sky130_fd_sc_hd__nand2_1 c512 (.A(net429),
    .B(net328),
    .Y(net435));
 sky130_fd_sc_hd__nor2_1 c513 (.A(net198),
    .B(net431),
    .Y(net436));
 sky130_fd_sc_hd__nand2_1 c514 (.A(net76),
    .B(net335),
    .Y(net437));
 sky130_fd_sc_hd__and2b_1 c515 (.A_N(net329),
    .B(net785),
    .X(net438));
 sky130_fd_sc_hd__nor2b_2 c516 (.A(net435),
    .B_N(net431),
    .Y(net439));
 sky130_fd_sc_hd__and2b_1 c517 (.A_N(net437),
    .B(net433),
    .X(net440));
 sky130_fd_sc_hd__dfrbp_1 c518 (.CLK(clknet_4_10_0_clk),
    .D(net429),
    .RESET_B(net440),
    .Q(net441));
 sky130_fd_sc_hd__nand2b_1 c519 (.A_N(net325),
    .B(net437),
    .Y(net442));
 sky130_fd_sc_hd__a21boi_2 c52 (.A1(net690),
    .A2(net712),
    .B1_N(net773),
    .Y(net0));
 sky130_fd_sc_hd__nand2b_1 c520 (.A_N(net435),
    .B(net433),
    .Y(net443));
 sky130_fd_sc_hd__nor2b_2 c521 (.A(net436),
    .B_N(net212),
    .Y(net444));
 sky130_fd_sc_hd__dfrtn_1 c522 (.CLK_N(clknet_4_10_0_clk),
    .D(net434),
    .RESET_B(net439),
    .Q(net445));
 sky130_fd_sc_hd__or2b_1 c523 (.A(net442),
    .B_N(net444),
    .X(net446));
 sky130_fd_sc_hd__or2b_2 c524 (.A(net444),
    .B_N(net436),
    .X(net447));
 sky130_fd_sc_hd__and2b_1 c525 (.A_N(net689),
    .B(net343),
    .X(net448));
 sky130_fd_sc_hd__o31a_1 c526 (.A1(net701),
    .A2(net431),
    .A3(net360),
    .B1(net326),
    .X(net449));
 sky130_fd_sc_hd__and2b_1 c527 (.A_N(net111),
    .B(net337),
    .X(net450));
 sky130_fd_sc_hd__dfrtp_1 c528 (.CLK(clknet_4_10_0_clk),
    .D(net216),
    .RESET_B(net439),
    .Q(net451));
 sky130_fd_sc_hd__nor2_1 c529 (.A(net450),
    .B(net793),
    .Y(net452));
 sky130_fd_sc_hd__a21oi_2 c53 (.A1(net710),
    .A2(net683),
    .B1(net713),
    .Y(net1));
 sky130_fd_sc_hd__dfrtp_1 c530 (.CLK(clknet_4_10_0_clk),
    .D(net443),
    .RESET_B(net445),
    .Q(net453));
 sky130_fd_sc_hd__nand2b_1 c531 (.A_N(net326),
    .B(net782),
    .Y(net454));
 sky130_fd_sc_hd__dfrtp_1 c532 (.CLK(clknet_4_10_0_clk),
    .D(net806),
    .RESET_B(net428),
    .Q(net455));
 sky130_fd_sc_hd__sdfxtp_1 c533 (.CLK(clknet_4_10_0_clk),
    .D(net428),
    .SCD(net443),
    .SCE(net344),
    .Q(net456));
 sky130_fd_sc_hd__or2_1 c534 (.A(net441),
    .B(net456),
    .X(net457));
 sky130_fd_sc_hd__or2_2 c535 (.A(net793),
    .B(net344),
    .X(net458));
 sky130_fd_sc_hd__dfsbp_1 c536 (.CLK(clknet_4_8_0_clk),
    .D(net452),
    .SET_B(net799),
    .Q(net459));
 sky130_fd_sc_hd__o31ai_1 c537 (.A1(net449),
    .A2(net455),
    .A3(net344),
    .B1(net444),
    .Y(net460));
 sky130_fd_sc_hd__a21oi_1 c538 (.A1(net232),
    .A2(net354),
    .B1(net449),
    .Y(net461));
 sky130_fd_sc_hd__o21ai_1 c539 (.A1(net431),
    .A2(net74),
    .B1(net714),
    .Y(net462));
 sky130_fd_sc_hd__o41a_2 c54 (.A1(net0),
    .A2(net705),
    .A3(net1),
    .A4(net704),
    .B1(net773),
    .X(net2));
 sky130_fd_sc_hd__a21o_1 c540 (.A1(net354),
    .A2(net460),
    .B1(net458),
    .X(net463));
 sky130_fd_sc_hd__o21a_2 c541 (.A1(net337),
    .A2(net209),
    .B1(net701),
    .X(net464));
 sky130_fd_sc_hd__nor2b_1 c542 (.A(net454),
    .B_N(net457),
    .Y(net465));
 sky130_fd_sc_hd__and2_4 c543 (.A(net459),
    .B(net464),
    .X(net737));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net432),
    .A1(net456),
    .A2(net461),
    .A3(net352),
    .S0(net737),
    .S1(net433),
    .X(net466));
 sky130_fd_sc_hd__sdfbbp_1 c545 (.CLK(clknet_4_10_0_clk),
    .D(net448),
    .RESET_B(net804),
    .SCD(net737),
    .SCE(net783),
    .SET_B(net344),
    .Q(net468),
    .Q_N(net467));
 sky130_fd_sc_hd__nor2_4 c546 (.A(net714),
    .B(clknet_1_1__leaf_net384),
    .Y(net469));
 sky130_fd_sc_hd__or2b_1 c547 (.A(net124),
    .B_N(net444),
    .X(net470));
 sky130_fd_sc_hd__and2b_1 c548 (.A_N(net122),
    .B(net242),
    .X(net471));
 sky130_fd_sc_hd__and2_0 c549 (.A(net242),
    .B(net470),
    .X(net472));
 sky130_fd_sc_hd__a21o_1 c55 (.A1(net707),
    .A2(net703),
    .B1(net708),
    .X(net3));
 sky130_fd_sc_hd__dfsbp_2 c550 (.CLK(clknet_4_14_0_clk),
    .D(net469),
    .SET_B(net737),
    .Q(net474),
    .Q_N(net473));
 sky130_fd_sc_hd__nor2_1 c551 (.A(net103),
    .B(net472),
    .Y(net475));
 sky130_fd_sc_hd__nor2_1 c552 (.A(net343),
    .B(net458),
    .Y(net476));
 sky130_fd_sc_hd__a21boi_1 c553 (.A1(net476),
    .A2(net127),
    .B1_N(clknet_1_1__leaf_net371),
    .Y(net477));
 sky130_fd_sc_hd__nand2_1 c554 (.A(net361),
    .B(net714),
    .Y(net478));
 sky130_fd_sc_hd__a21oi_1 c555 (.A1(net355),
    .A2(net474),
    .B1(net458),
    .Y(net479));
 sky130_fd_sc_hd__and2b_1 c556 (.A_N(net465),
    .B(net363),
    .X(net480));
 sky130_fd_sc_hd__mux4_4 c557 (.A0(net332),
    .A1(net477),
    .A2(clknet_1_0__leaf_net377),
    .A3(net737),
    .S0(net479),
    .S1(net343),
    .X(net481));
 sky130_fd_sc_hd__dfstp_1 c558 (.CLK(clknet_4_12_0_clk),
    .D(net475),
    .SET_B(net127),
    .Q(net482));
 sky130_fd_sc_hd__dfbbn_1 c559 (.CLK_N(clknet_4_9_0_clk),
    .D(net479),
    .RESET_B(net252),
    .SET_B(net471),
    .Q(net483));
 sky130_fd_sc_hd__o41a_1 c56 (.A1(net696),
    .A2(net3),
    .A3(net706),
    .A4(net698),
    .B1(net773),
    .X(net4));
 sky130_fd_sc_hd__nor2b_1 c560 (.A(net367),
    .B_N(net474),
    .Y(net484));
 sky130_fd_sc_hd__sdfstp_1 c561 (.CLK(clknet_4_9_0_clk),
    .D(net372),
    .SCD(clknet_1_0__leaf_net381),
    .SCE(clknet_1_0__leaf_net384),
    .SET_B(net737),
    .Q(net485));
 sky130_fd_sc_hd__o31ai_4 c562 (.A1(clknet_1_1__leaf_net371),
    .A2(net367),
    .A3(net485),
    .B1(net473),
    .Y(net486));
 sky130_fd_sc_hd__dfstp_1 c563 (.CLK(clknet_4_12_0_clk),
    .D(net378),
    .SET_B(net803),
    .Q(net487));
 sky130_fd_sc_hd__nor2b_2 c564 (.A(net485),
    .B_N(net487),
    .Y(net488));
 sky130_fd_sc_hd__o41a_4 c565 (.A1(net480),
    .A2(clknet_1_0__leaf_net486),
    .A3(net444),
    .A4(net487),
    .B1(net465),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net471),
    .A1(clknet_1_0__leaf_net489),
    .A2(net343),
    .A3(net132),
    .S0(clknet_1_1__leaf_net486),
    .S1(net656),
    .X(net490));
 sky130_fd_sc_hd__mux2_8 c567 (.A0(net28),
    .A1(net93),
    .S(clknet_1_1__leaf_net381),
    .X(net491));
 sky130_fd_sc_hd__dfstp_1 c568 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net491),
    .SET_B(net737),
    .Q(net492));
 sky130_fd_sc_hd__dfbbn_1 c569 (.CLK_N(clknet_4_12_0_clk),
    .D(net682),
    .RESET_B(net252),
    .SET_B(net492),
    .Q(net493));
 sky130_fd_sc_hd__o21ai_4 c57 (.A1(net708),
    .A2(net712),
    .B1(net2),
    .Y(net5));
 sky130_fd_sc_hd__dfbbp_1 c570 (.CLK(clknet_4_12_0_clk),
    .D(net440),
    .RESET_B(net458),
    .SET_B(clknet_1_0__leaf_net491),
    .Q(net495),
    .Q_N(net494));
 sky130_fd_sc_hd__and2_1 c571 (.A(net478),
    .B(net492),
    .X(net496));
 sky130_fd_sc_hd__a21boi_4 c572 (.A1(clknet_1_0__leaf_net389),
    .A2(clknet_1_0__leaf_net491),
    .B1_N(net392),
    .Y(net497));
 sky130_fd_sc_hd__sdfxbp_1 c573 (.CLK(clknet_4_12_0_clk),
    .D(net375),
    .SCD(net493),
    .SCE(net492),
    .Q(net498));
 sky130_fd_sc_hd__o21ba_2 c574 (.A1(net492),
    .A2(net339),
    .B1_N(clknet_1_1__leaf_net389),
    .X(net499));
 sky130_fd_sc_hd__mux4_2 c575 (.A0(net496),
    .A1(net24),
    .A2(clknet_1_1__leaf_net491),
    .A3(clknet_1_1__leaf_net388),
    .S0(net729),
    .S1(net494),
    .X(net500));
 sky130_fd_sc_hd__dlrbn_2 c576 (.D(clknet_1_1__leaf_net381),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net405),
    .Q(net763),
    .Q_N(net501));
 sky130_fd_sc_hd__dlrbn_1 c577 (.D(net497),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net499),
    .Q(net503),
    .Q_N(net502));
 sky130_fd_sc_hd__o21ai_0 c578 (.A1(net498),
    .A2(net740),
    .B1(net501),
    .Y(net504));
 sky130_fd_sc_hd__or2b_1 c579 (.A(net784),
    .B_N(net502),
    .X(net505));
 sky130_fd_sc_hd__o31ai_1 c58 (.A1(net4),
    .A2(net680),
    .A3(net690),
    .B1(net773),
    .Y(net6));
 sky130_fd_sc_hd__and2b_1 c580 (.A_N(net505),
    .B(net763),
    .X(net506));
 sky130_fd_sc_hd__o31ai_1 c581 (.A1(net135),
    .A2(net506),
    .A3(clknet_1_1__leaf_net381),
    .B1(net501),
    .Y(net507));
 sky130_fd_sc_hd__or2b_1 c582 (.A(net339),
    .B_N(net503),
    .X(net508));
 sky130_fd_sc_hd__nand2b_2 c583 (.A_N(net504),
    .B(net506),
    .Y(net509));
 sky130_fd_sc_hd__nand2b_1 c584 (.A_N(clknet_1_0__leaf_net507),
    .B(net470),
    .Y(net510));
 sky130_fd_sc_hd__sdfxbp_1 c585 (.CLK(clknet_4_13_0_clk),
    .D(net508),
    .SCD(net510),
    .SCE(net458),
    .Q(net511));
 sky130_fd_sc_hd__or2_1 c586 (.A(net383),
    .B(net509),
    .X(net512));
 sky130_fd_sc_hd__mux4_2 c587 (.A0(net512),
    .A1(net511),
    .A2(clknet_1_1__leaf_net507),
    .A3(net509),
    .S0(net382),
    .S1(net494),
    .X(net513));
 sky130_fd_sc_hd__o21ai_1 c588 (.A1(net503),
    .A2(net363),
    .B1(net671),
    .Y(net514));
 sky130_fd_sc_hd__or2_1 c589 (.A(net407),
    .B(net509),
    .X(net515));
 sky130_fd_sc_hd__a21o_1 c59 (.A1(net703),
    .A2(net706),
    .B1(net6),
    .X(net7));
 sky130_fd_sc_hd__o21ba_1 c590 (.A1(net487),
    .A2(net506),
    .B1_N(net742),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 c591 (.A(net664),
    .X(net517));
 sky130_fd_sc_hd__a21o_1 c592 (.A1(net155),
    .A2(net421),
    .B1(net744),
    .X(net518));
 sky130_fd_sc_hd__o21ai_1 c593 (.A1(net141),
    .A2(net763),
    .B1(net740),
    .Y(net519));
 sky130_fd_sc_hd__a21bo_1 c594 (.A1(net482),
    .A2(net339),
    .B1_N(net458),
    .X(net520));
 sky130_fd_sc_hd__a21o_2 c595 (.A1(net392),
    .A2(clknet_1_0__leaf_net749),
    .B1(net509),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_2 c596 (.A(net805),
    .X(net736));
 sky130_fd_sc_hd__mux4_2 c597 (.A0(net166),
    .A1(net517),
    .A2(net506),
    .A3(net736),
    .S0(clknet_1_0__leaf_net749),
    .S1(net407),
    .X(net522));
 sky130_fd_sc_hd__sdfstp_1 c598 (.CLK(clknet_4_13_0_clk),
    .D(net520),
    .SCD(net474),
    .SCE(clknet_1_0__leaf_net513),
    .SET_B(net736),
    .Q(net523));
 sky130_fd_sc_hd__mux4_4 c599 (.A0(net519),
    .A1(net171),
    .A2(net676),
    .A3(net736),
    .S0(net473),
    .S1(net517),
    .X(net524));
 sky130_fd_sc_hd__o21ai_4 c60 (.A1(net5),
    .A2(net701),
    .B1(net680),
    .Y(net8));
 sky130_fd_sc_hd__o31a_1 c600 (.A1(net281),
    .A2(clknet_1_0__leaf_net388),
    .A3(clknet_1_0__leaf_net750),
    .B1(net657),
    .X(net525));
 sky130_fd_sc_hd__o21ba_1 c601 (.A1(net446),
    .A2(net474),
    .B1_N(net658),
    .X(net526));
 sky130_fd_sc_hd__sdfxtp_1 c602 (.CLK(clknet_4_13_0_clk),
    .D(net252),
    .SCD(net525),
    .SCE(net676),
    .Q(net527));
 sky130_fd_sc_hd__sdfxtp_1 c603 (.CLK(clknet_4_13_0_clk),
    .D(net518),
    .SCD(net736),
    .SCE(net509),
    .Q(net528));
 sky130_fd_sc_hd__sdfstp_1 c604 (.CLK(clknet_4_13_0_clk),
    .D(net809),
    .SCD(net526),
    .SCE(net737),
    .SET_B(net838),
    .Q(net748));
 sky130_fd_sc_hd__sdfxtp_1 c605 (.CLK(clknet_4_13_0_clk),
    .D(net363),
    .SCD(clknet_1_0__leaf_net513),
    .SCE(net204),
    .Q(net529));
 sky130_fd_sc_hd__sdfbbn_1 c606 (.CLK_N(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net500),
    .RESET_B(net736),
    .SCD(clknet_1_1__leaf_net513),
    .SCE(net526),
    .SET_B(net171),
    .Q(net530));
 sky130_fd_sc_hd__a21boi_1 c607 (.A1(net528),
    .A2(net458),
    .B1_N(net740),
    .Y(net531));
 sky130_fd_sc_hd__a21o_1 c608 (.A1(net495),
    .A2(net529),
    .B1(net531),
    .X(net532));
 sky130_fd_sc_hd__o21ba_1 c61 (.A1(net680),
    .A2(net7),
    .B1_N(net4),
    .X(net9));
 sky130_fd_sc_hd__o21ai_1 c62 (.A1(net8),
    .A2(net9),
    .B1(net678),
    .Y(net10));
 sky130_fd_sc_hd__or2_2 c63 (.A(net698),
    .B(net12),
    .X(net11));
 sky130_fd_sc_hd__and2b_1 c630 (.A_N(net324),
    .B(net751),
    .X(net533));
 sky130_fd_sc_hd__and2_1 c631 (.A(net438),
    .B(net445),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_1 c632 (.A(net637),
    .X(net535));
 sky130_fd_sc_hd__inv_2 c633 (.A(net637),
    .Y(net536));
 sky130_fd_sc_hd__dlrbp_1 c634 (.D(net439),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net204),
    .Q(net538),
    .Q_N(net537));
 sky130_fd_sc_hd__nand2_1 c635 (.A(net711),
    .B(net534),
    .Y(net539));
 sky130_fd_sc_hd__and2b_1 c636 (.A_N(net676),
    .B(net445),
    .X(net540));
 sky130_fd_sc_hd__nor2_2 c637 (.A(net679),
    .B(net537),
    .Y(net541));
 sky130_fd_sc_hd__dlrbp_1 c638 (.D(net785),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net434),
    .Q(net543),
    .Q_N(net542));
 sky130_fd_sc_hd__nand2b_1 c639 (.A_N(net534),
    .B(net751),
    .Y(net544));
 sky130_fd_sc_hd__nor2b_4 c64 (.A(net707),
    .B_N(net5),
    .Y(net721));
 sky130_fd_sc_hd__or2_1 c640 (.A(net535),
    .B(net542),
    .X(net545));
 sky130_fd_sc_hd__nand2b_2 c641 (.A_N(net543),
    .B(net679),
    .Y(net546));
 sky130_fd_sc_hd__dlrtn_1 c642 (.D(net334),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net534),
    .Q(net547));
 sky130_fd_sc_hd__dlrtn_1 c643 (.D(net338),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net209),
    .Q(net548));
 sky130_fd_sc_hd__nor2b_1 c644 (.A(net548),
    .B_N(net541),
    .Y(net549));
 sky130_fd_sc_hd__and2_1 c645 (.A(net547),
    .B(net539),
    .X(net550));
 sky130_fd_sc_hd__dlrtn_2 c646 (.D(net544),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net825),
    .Q(net551));
 sky130_fd_sc_hd__o21ba_1 c647 (.A1(net550),
    .A2(net551),
    .B1_N(net537),
    .X(net552));
 sky130_fd_sc_hd__dlrtp_1 c648 (.D(net552),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net538),
    .Q(net553));
 sky130_fd_sc_hd__a21o_1 c649 (.A1(net553),
    .A2(net438),
    .B1(net816),
    .X(net554));
 sky130_fd_sc_hd__and2_2 c65 (.A(net673),
    .B(net715),
    .X(net12));
 sky130_fd_sc_hd__dfbbn_1 c650 (.CLK_N(clknet_4_10_0_clk),
    .D(net534),
    .RESET_B(net554),
    .SET_B(net552),
    .Q(net556),
    .Q_N(net555));
 sky130_fd_sc_hd__and2_2 c651 (.A(net461),
    .B(net672),
    .X(net557));
 sky130_fd_sc_hd__and2_2 c652 (.A(net113),
    .B(net538),
    .X(net558));
 sky130_fd_sc_hd__dlrtp_1 c653 (.D(net540),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net557),
    .Q(net559));
 sky130_fd_sc_hd__o41a_1 c654 (.A1(net457),
    .A2(net781),
    .A3(net558),
    .A4(net468),
    .B1(net541),
    .X(net560));
 sky130_fd_sc_hd__nand2_1 c655 (.A(net558),
    .B(net93),
    .Y(net561));
 sky130_fd_sc_hd__mux4_1 c656 (.A0(net352),
    .A1(net468),
    .A2(net555),
    .A3(net711),
    .S0(net558),
    .S1(net557),
    .X(net562));
 sky130_fd_sc_hd__or2_2 c657 (.A(net238),
    .B(net540),
    .X(net563));
 sky130_fd_sc_hd__dlrtp_2 c658 (.D(net462),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net557),
    .Q(net564));
 sky130_fd_sc_hd__edfxbp_1 c659 (.CLK(clknet_4_11_0_clk),
    .D(net557),
    .DE(net546),
    .Q(net565));
 sky130_fd_sc_hd__or2b_1 c66 (.A(net6),
    .B_N(net707),
    .X(net13));
 sky130_fd_sc_hd__or2b_1 c660 (.A(net463),
    .B_N(net558),
    .X(net566));
 sky130_fd_sc_hd__and2_1 c661 (.A(net565),
    .B(net462),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c662 (.A0(net561),
    .A1(net209),
    .A2(net751),
    .A3(net557),
    .S0(net563),
    .S1(net238),
    .X(net568));
 sky130_fd_sc_hd__or2_1 c663 (.A(net468),
    .B(net564),
    .X(net569));
 sky130_fd_sc_hd__and2b_2 c664 (.A_N(net566),
    .B(net564),
    .X(net570));
 sky130_fd_sc_hd__and2_0 c665 (.A(net556),
    .B(net655),
    .X(net571));
 sky130_fd_sc_hd__and2_1 c666 (.A(net560),
    .B(net571),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(net347),
    .A1(net751),
    .A2(net557),
    .A3(net734),
    .S0(net570),
    .S1(net549),
    .X(net573));
 sky130_fd_sc_hd__o21ai_1 c668 (.A1(net570),
    .A2(net467),
    .B1(net659),
    .Y(net574));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_4_11_0_clk),
    .D(net439),
    .RESET_B(net558),
    .SCD(net467),
    .SCE(net464),
    .SET_B(net661),
    .Q(net575));
 sky130_fd_sc_hd__or2_2 c67 (.A(net674),
    .B(net5),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net464),
    .A1(net558),
    .A2(net541),
    .A3(net536),
    .S0(net433),
    .S1(net832),
    .X(net576));
 sky130_fd_sc_hd__edfxtp_1 c671 (.CLK(clknet_4_11_0_clk),
    .D(net576),
    .DE(net575),
    .Q(net577));
 sky130_fd_sc_hd__nor2_1 c672 (.A(net445),
    .B(net549),
    .Y(net578));
 sky130_fd_sc_hd__or2b_2 c673 (.A(net569),
    .B_N(net537),
    .X(net725));
 sky130_fd_sc_hd__nand2b_1 c674 (.A_N(net572),
    .B(net751),
    .Y(net579));
 sky130_fd_sc_hd__and2b_1 c675 (.A_N(net559),
    .B(net570),
    .X(net580));
 sky130_fd_sc_hd__o41a_4 c676 (.A1(net538),
    .A2(clknet_1_0__leaf_net489),
    .A3(net751),
    .A4(net577),
    .B1(net563),
    .X(net581));
 sky130_fd_sc_hd__dfbbn_1 c677 (.CLK_N(clknet_4_15_0_clk),
    .D(clknet_1_0__leaf_net377),
    .RESET_B(clknet_1_1__leaf_net581),
    .SET_B(net672),
    .Q(net582));
 sky130_fd_sc_hd__dfbbp_1 c678 (.CLK(clknet_4_11_0_clk),
    .D(net483),
    .RESET_B(clknet_1_0__leaf_net581),
    .SET_B(net577),
    .Q(net584),
    .Q_N(net583));
 sky130_fd_sc_hd__a21oi_1 c679 (.A1(net132),
    .A2(net551),
    .B1(net541),
    .Y(net585));
 sky130_fd_sc_hd__nor2_1 c68 (.A(net13),
    .B(net1),
    .Y(net15));
 sky130_fd_sc_hd__sedfxbp_1 c680 (.CLK(clknet_4_15_0_clk),
    .D(net582),
    .DE(clknet_1_1__leaf_net581),
    .SCD(clknet_1_1__leaf_net489),
    .SCE(clknet_1_1__leaf_net377),
    .Q(net586));
 sky130_fd_sc_hd__sdfxbp_1 c681 (.CLK(clknet_4_14_0_clk),
    .D(net578),
    .SCD(net464),
    .SCE(clknet_1_0__leaf_net581),
    .Q(net587));
 sky130_fd_sc_hd__inv_1 c682 (.A(net835),
    .Y(net588));
 sky130_fd_sc_hd__inv_6 c683 (.A(net641),
    .Y(net589));
 sky130_fd_sc_hd__o21ai_2 c684 (.A1(net545),
    .A2(net588),
    .B1(net577),
    .Y(net590));
 sky130_fd_sc_hd__sdfxbp_1 c685 (.CLK(clknet_4_11_0_clk),
    .D(net580),
    .SCD(net590),
    .SCE(net588),
    .Q(net592),
    .Q_N(net591));
 sky130_fd_sc_hd__sdfxtp_1 c686 (.CLK(clknet_4_14_0_clk),
    .D(net585),
    .SCD(net821),
    .SCE(net580),
    .Q(net593));
 sky130_fd_sc_hd__o41a_1 c687 (.A1(net127),
    .A2(net593),
    .A3(net725),
    .A4(net590),
    .B1(net584),
    .X(net594));
 sky130_fd_sc_hd__o41a_1 c688 (.A1(net567),
    .A2(net589),
    .A3(net445),
    .A4(net577),
    .B1(net488),
    .X(net595));
 sky130_fd_sc_hd__o21bai_4 c689 (.A1(net551),
    .A2(net589),
    .B1_N(net595),
    .Y(net722));
 sky130_fd_sc_hd__and2_1 c69 (.A(net678),
    .B(net843),
    .X(net16));
 sky130_fd_sc_hd__o31a_1 c690 (.A1(net484),
    .A2(net595),
    .A3(net722),
    .B1(net594),
    .X(net596));
 sky130_fd_sc_hd__o41a_2 c691 (.A1(clknet_1_1__leaf_net384),
    .A2(net595),
    .A3(net464),
    .A4(net591),
    .B1(net563),
    .X(net597));
 sky130_fd_sc_hd__mux2_1 c692 (.A0(net594),
    .A1(net722),
    .S(net595),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_1 c693 (.A(net663),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_1 c694 (.A(net663),
    .X(net599));
 sky130_fd_sc_hd__sdfxtp_1 c695 (.CLK(clknet_4_14_0_clk),
    .D(net830),
    .SCD(net277),
    .SCE(net729),
    .Q(net719));
 sky130_fd_sc_hd__o21bai_1 c696 (.A1(net563),
    .A2(net145),
    .B1_N(net734),
    .Y(net600));
 sky130_fd_sc_hd__o21a_1 c697 (.A1(net433),
    .A2(net771),
    .B1(net702),
    .X(net601));
 sky130_fd_sc_hd__sdfxtp_1 c698 (.CLK(clknet_4_14_0_clk),
    .D(net601),
    .SCD(net779),
    .SCE(net495),
    .Q(net602));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net570),
    .A1(net592),
    .A2(net433),
    .A3(net725),
    .S0(net494),
    .S1(net577),
    .X(net603));
 sky130_fd_sc_hd__and2_1 c70 (.A(net843),
    .B(net11),
    .X(net17));
 sky130_fd_sc_hd__a21o_1 c700 (.A1(net536),
    .A2(net672),
    .B1(net570),
    .X(net604));
 sky130_fd_sc_hd__dfbbn_1 c701 (.CLK_N(clknet_4_11_0_clk),
    .D(net79),
    .RESET_B(net604),
    .SET_B(net564),
    .Q(net605));
 sky130_fd_sc_hd__or2b_1 c702 (.A(net464),
    .B_N(net596),
    .X(net606));
 sky130_fd_sc_hd__dfbbn_1 c703 (.CLK_N(clknet_4_15_0_clk),
    .D(net606),
    .RESET_B(net495),
    .SET_B(net823),
    .Q(net608),
    .Q_N(net607));
 sky130_fd_sc_hd__dfbbp_1 c704 (.CLK(clknet_4_14_0_clk),
    .D(net277),
    .RESET_B(net577),
    .SET_B(net601),
    .Q(net610),
    .Q_N(net609));
 sky130_fd_sc_hd__and2_0 c705 (.A(net610),
    .B(net495),
    .X(net611));
 sky130_fd_sc_hd__a21o_1 c706 (.A1(net587),
    .A2(net21),
    .B1(net607),
    .X(net612));
 sky130_fd_sc_hd__mux4_4 c707 (.A0(net600),
    .A1(net145),
    .A2(net609),
    .A3(net591),
    .S0(net501),
    .S1(net570),
    .X(net613));
 sky130_fd_sc_hd__mux2_1 c708 (.A0(net24),
    .A1(net605),
    .S(net564),
    .X(net614));
 sky130_fd_sc_hd__a21o_1 c709 (.A1(net541),
    .A2(net599),
    .B1(net209),
    .X(net727));
 sky130_fd_sc_hd__nor2_1 c71 (.A(net11),
    .B(net677),
    .Y(net18));
 sky130_fd_sc_hd__mux2_1 c710 (.A0(net612),
    .A1(net611),
    .S(net464),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net613),
    .A1(net574),
    .A2(net546),
    .A3(clknet_1_0__leaf_net489),
    .S0(net564),
    .S1(net596),
    .X(net616));
 sky130_fd_sc_hd__a21oi_1 c712 (.A1(net614),
    .A2(net584),
    .B1(net662),
    .Y(net617));
 sky130_fd_sc_hd__sdfxbp_1 c713 (.CLK(clknet_4_15_0_clk),
    .D(net608),
    .SCD(net671),
    .SCE(clknet_1_1__leaf_net581),
    .Q(net618));
 sky130_fd_sc_hd__a21bo_1 c714 (.A1(net516),
    .A2(net93),
    .B1_N(net729),
    .X(net619));
 sky130_fd_sc_hd__inv_6 c715 (.A(net635),
    .Y(net726));
 sky130_fd_sc_hd__sedfxbp_1 c716 (.CLK(clknet_4_15_0_clk),
    .D(net549),
    .DE(net615),
    .SCD(clknet_1_1__leaf_net489),
    .SCE(net546),
    .Q(net620));
 sky130_fd_sc_hd__o41a_1 c717 (.A1(net209),
    .A2(net530),
    .A3(net598),
    .A4(net93),
    .B1(net778),
    .X(net621));
 sky130_fd_sc_hd__o31a_1 c718 (.A1(net488),
    .A2(net523),
    .A3(clknet_1_1__leaf_net388),
    .B1(net204),
    .X(net622));
 sky130_fd_sc_hd__mux2_8 c719 (.A0(net602),
    .A1(clknet_1_1__leaf_net489),
    .S(net734),
    .X(net623));
 sky130_fd_sc_hd__a21boi_2 c72 (.A1(net683),
    .A2(net18),
    .B1_N(net721),
    .Y(net19));
 sky130_fd_sc_hd__o21a_1 c720 (.A1(net447),
    .A2(net619),
    .B1(net722),
    .X(net624));
 sky130_fd_sc_hd__inv_1 c721 (.A(net635),
    .Y(net625));
 sky130_fd_sc_hd__sedfxtp_2 c722 (.CLK(clknet_4_15_0_clk),
    .D(net93),
    .DE(net590),
    .SCD(net447),
    .SCE(net424),
    .Q(net626));
 sky130_fd_sc_hd__o31a_1 c723 (.A1(net620),
    .A2(net626),
    .A3(net488),
    .B1(net657),
    .X(net627));
 sky130_fd_sc_hd__sdfxbp_1 c724 (.CLK(clknet_4_15_0_clk),
    .D(net623),
    .SCD(net624),
    .SCE(net204),
    .Q(net628));
 sky130_fd_sc_hd__o21a_2 c725 (.A1(net546),
    .A2(net598),
    .B1(net626),
    .X(net629));
 sky130_fd_sc_hd__o21a_1 c726 (.A1(net628),
    .A2(net618),
    .B1(net702),
    .X(net630));
 sky130_fd_sc_hd__o41a_1 c727 (.A1(net627),
    .A2(net625),
    .A3(net771),
    .A4(net447),
    .B1(net501),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net586),
    .A1(net631),
    .A2(net629),
    .A3(net626),
    .S0(net719),
    .S1(net657),
    .X(net728));
 sky130_fd_sc_hd__sdfxtp_1 c729 (.CLK(clknet_4_15_0_clk),
    .D(clknet_1_1__leaf_net581),
    .SCD(net621),
    .SCE(net725),
    .Q(net720));
 sky130_fd_sc_hd__and2_1 c73 (.A(net19),
    .B(net16),
    .X(net20));
 sky130_fd_sc_hd__a21boi_4 c730 (.A1(net629),
    .A2(net622),
    .B1_N(net768),
    .Y(net632));
 sky130_fd_sc_hd__o21ai_1 c731 (.A1(net702),
    .A2(net532),
    .B1(net768),
    .Y(net633));
 sky130_fd_sc_hd__o31ai_1 c732 (.A1(net630),
    .A2(net515),
    .A3(net768),
    .B1(net626),
    .Y(net634));
 sky130_fd_sc_hd__o31ai_2 c733 (.A1(net633),
    .A2(net617),
    .A3(net447),
    .B1(net629),
    .Y(net741));
 sky130_fd_sc_hd__sdfxtp_2 c734 (.CLK(clknet_4_15_0_clk),
    .D(net634),
    .SCD(net632),
    .SCE(net629));
 sky130_fd_sc_hd__o21bai_4 c74 (.A1(net14),
    .A2(net17),
    .B1_N(net19),
    .Y(net21));
 sky130_fd_sc_hd__or2b_1 c75 (.A(net20),
    .B_N(net21),
    .X(net22));
 sky130_fd_sc_hd__and2_1 c76 (.A(net18),
    .B(net19),
    .X(net23));
 sky130_fd_sc_hd__mux2_2 c77 (.A0(net13),
    .A1(net699),
    .S(net698),
    .X(net24));
 sky130_fd_sc_hd__and2b_2 c78 (.A_N(net16),
    .B(net19),
    .X(net25));
 sky130_fd_sc_hd__nor2_1 c79 (.A(net25),
    .B(net15),
    .Y(net26));
 sky130_fd_sc_hd__o31ai_4 c80 (.A1(net705),
    .A2(net22),
    .A3(net26),
    .B1(net25),
    .Y(net27));
 sky130_fd_sc_hd__o31ai_4 c81 (.A1(net21),
    .A2(net27),
    .A3(net23),
    .B1(net678),
    .Y(net766));
 sky130_fd_sc_hd__o21ai_2 c82 (.A1(net26),
    .A2(net25),
    .B1(net20),
    .Y(net28));
 sky130_fd_sc_hd__o31ai_2 c83 (.A1(net22),
    .A2(net27),
    .A3(net21),
    .B1(net774),
    .Y(net29));
 sky130_fd_sc_hd__clkbuf_1 c84 (.A(net25),
    .X(net30));
 sky130_fd_sc_hd__inv_1 c85 (.A(net699),
    .Y(net31));
 sky130_fd_sc_hd__clkbuf_1 c86 (.A(net7),
    .X(net32));
 sky130_fd_sc_hd__or2b_1 c87 (.A(net30),
    .B_N(net32),
    .X(net33));
 sky130_fd_sc_hd__nand2_1 c88 (.A(net710),
    .B(net12),
    .Y(net34));
 sky130_fd_sc_hd__or2_1 c89 (.A(net30),
    .B(net11),
    .X(net35));
 sky130_fd_sc_hd__nor2_1 c90 (.A(net9),
    .B(net3),
    .Y(net36));
 sky130_fd_sc_hd__nand2_1 c91 (.A(net35),
    .B(net30),
    .Y(net37));
 sky130_fd_sc_hd__and2_1 c92 (.A(net34),
    .B(net36),
    .X(net38));
 sky130_fd_sc_hd__and2_1 c93 (.A(net35),
    .B(net34),
    .X(net39));
 sky130_fd_sc_hd__o21bai_2 c94 (.A1(net3),
    .A2(net36),
    .B1_N(net12),
    .Y(net40));
 sky130_fd_sc_hd__nand2b_1 c95 (.A_N(net40),
    .B(net36),
    .Y(net41));
 sky130_fd_sc_hd__nor2_1 c96 (.A(net36),
    .B(net38),
    .Y(net42));
 sky130_fd_sc_hd__or2_2 c97 (.A(net37),
    .B(net39),
    .X(net43));
 sky130_fd_sc_hd__nor2_1 c98 (.A(net43),
    .B(net15),
    .Y(net44));
 sky130_fd_sc_hd__nand2b_2 c99 (.A_N(net44),
    .B(net14),
    .Y(net45));
 sky130_fd_sc_hd__sedfxtp_4 merge755 (.CLK(clknet_4_15_0_clk),
    .D(net539),
    .DE(net603),
    .SCD(net424),
    .SCE(clknet_1_1__leaf_net388),
    .Q(net635));
 sky130_fd_sc_hd__mux4_4 merge756 (.A0(net117),
    .A1(net597),
    .A2(net464),
    .A3(net583),
    .S0(net494),
    .S1(clknet_1_0__leaf_net581),
    .X(net636));
 sky130_fd_sc_hd__sedfxtp_1 merge757 (.CLK(clknet_4_10_0_clk),
    .D(net74),
    .DE(net439),
    .SCD(net533),
    .SCE(net433),
    .Q(net637));
 sky130_fd_sc_hd__sdfrbp_1 merge758 (.CLK(clknet_4_6_0_clk),
    .D(net152),
    .RESET_B(net40),
    .SCD(net44),
    .SCE(net157),
    .Q(net639),
    .Q_N(net638));
 sky130_fd_sc_hd__mux4_2 merge759 (.A0(net514),
    .A1(net473),
    .A2(clknet_1_0__leaf_net500),
    .A3(net521),
    .S0(net744),
    .S1(net166),
    .X(net640));
 sky130_fd_sc_hd__sdfrbp_1 merge760 (.CLK(clknet_4_11_0_clk),
    .D(net579),
    .RESET_B(net132),
    .SCD(net490),
    .SCE(net580),
    .Q(net642),
    .Q_N(net641));
 sky130_fd_sc_hd__mux4_1 merge761 (.A0(net114),
    .A1(net302),
    .A2(net141),
    .A3(net290),
    .S0(net171),
    .S1(net771),
    .X(net643));
 sky130_fd_sc_hd__dfxbp_1 s762 (.CLK(clknet_4_5_0_clk),
    .D(net173),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__dfxbp_1 s763 (.CLK(clknet_4_5_0_clk),
    .D(net187),
    .Q(net646));
 sky130_fd_sc_hd__dfxtp_1 s764 (.CLK(clknet_4_5_0_clk),
    .D(net193),
    .Q(net647));
 sky130_fd_sc_hd__dfxtp_1 s765 (.CLK(clknet_4_6_0_clk),
    .D(net253),
    .Q(net648));
 sky130_fd_sc_hd__dfxtp_1 s766 (.CLK(clknet_4_9_0_clk),
    .D(net257),
    .Q(net649));
 sky130_fd_sc_hd__dlclkp_1 s767 (.CLK(clknet_4_6_0_clk),
    .GATE(net268),
    .GCLK(net650));
 sky130_fd_sc_hd__dlclkp_2 s768 (.CLK(clknet_4_7_0_clk),
    .GATE(net278),
    .GCLK(net651));
 sky130_fd_sc_hd__dlclkp_4 s769 (.CLK(clknet_4_3_0_clk),
    .GATE(net415),
    .GCLK(net652));
 sky130_fd_sc_hd__dlxbn_1 s770 (.D(net422),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net653));
 sky130_fd_sc_hd__dlxbn_1 s771 (.D(net423),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net654));
 sky130_fd_sc_hd__dlxbp_1 s772 (.D(net466),
    .GATE(clknet_4_10_0_clk),
    .Q(net655));
 sky130_fd_sc_hd__dlxtn_1 s773 (.D(net481),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net656));
 sky130_fd_sc_hd__dlxtn_1 s774 (.D(net522),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net657));
 sky130_fd_sc_hd__dlxtn_1 s775 (.D(net524),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net658));
 sky130_fd_sc_hd__dlxtp_1 s776 (.D(net562),
    .GATE(clknet_4_11_0_clk),
    .Q(net659));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s777 (.D(net568),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net660));
 sky130_fd_sc_hd__dfxbp_1 s778 (.CLK(clknet_4_11_0_clk),
    .D(net573),
    .Q(net661));
 sky130_fd_sc_hd__dfxbp_1 s779 (.CLK(clknet_4_14_0_clk),
    .D(net616),
    .Q(net662));
 sky130_fd_sc_hd__dfxtp_1 s780 (.CLK(clknet_4_14_0_clk),
    .D(net636),
    .Q(net663));
 sky130_fd_sc_hd__dfxtp_1 s781 (.CLK(clknet_4_3_0_clk),
    .D(net640),
    .Q(net664));
 sky130_fd_sc_hd__dfxtp_1 s782 (.CLK(clknet_4_3_0_clk),
    .D(net643),
    .Q(net665));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net667));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net668));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net669));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net670));
 sky130_fd_sc_hd__buf_6 input6 (.A(in13),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(in14),
    .X(net672));
 sky130_fd_sc_hd__buf_2 input8 (.A(in15),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net674));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net675));
 sky130_fd_sc_hd__buf_2 input11 (.A(in18),
    .X(net676));
 sky130_fd_sc_hd__buf_2 input12 (.A(in19),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(in2),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net679));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(in21),
    .X(net680));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net681));
 sky130_fd_sc_hd__buf_2 input17 (.A(in23),
    .X(net682));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net683));
 sky130_fd_sc_hd__buf_1 input19 (.A(in25),
    .X(net684));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net687));
 sky130_fd_sc_hd__buf_1 input23 (.A(in29),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in3),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net690));
 sky130_fd_sc_hd__buf_1 input26 (.A(in31),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(in32),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(in33),
    .X(net693));
 sky130_fd_sc_hd__buf_1 input29 (.A(in34),
    .X(net694));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(in37),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(in38),
    .X(net698));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(in4),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(in40),
    .X(net701));
 sky130_fd_sc_hd__buf_2 input37 (.A(in41),
    .X(net702));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net703));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in44),
    .X(net705));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net706));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net707));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(in47),
    .X(net708));
 sky130_fd_sc_hd__buf_1 input44 (.A(in48),
    .X(net709));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net710));
 sky130_fd_sc_hd__buf_2 input46 (.A(in5),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(in50),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(in6),
    .X(net714));
 sky130_fd_sc_hd__buf_8 input50 (.A(in7),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(in8),
    .X(net716));
 sky130_fd_sc_hd__buf_1 input52 (.A(in9),
    .X(net717));
 sky130_fd_sc_hd__buf_2 output53 (.A(net718),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net719),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net720),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output56 (.A(net841),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output57 (.A(net722),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output58 (.A(net723),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output59 (.A(net724),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output60 (.A(net725),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net726),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net727),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net728),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net729),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output65 (.A(net730),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output66 (.A(net731),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output67 (.A(net732),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output68 (.A(net733),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net734),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output70 (.A(net735),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output71 (.A(net736),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net737),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net738),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output74 (.A(net739),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output75 (.A(net740),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net741),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output77 (.A(net742),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output78 (.A(net743),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output79 (.A(net744),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output80 (.A(net745),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output81 (.A(net746),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output82 (.A(net747),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output83 (.A(net748),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(clknet_1_1__leaf_net749),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(clknet_1_1__leaf_net750),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output86 (.A(net751),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output87 (.A(net777),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output88 (.A(net753),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output89 (.A(net754),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output90 (.A(net755),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output91 (.A(net756),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output92 (.A(net757),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output93 (.A(net758),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output94 (.A(net759),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output95 (.A(net760),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output96 (.A(net761),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output97 (.A(net762),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net763),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output99 (.A(net764),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output100 (.A(net765),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output101 (.A(net766),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net767),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output103 (.A(net768),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output104 (.A(net769),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(net225),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_2 max_cap106 (.A(net766),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(net743),
    .X(net772));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(net774),
    .X(net773));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(net713),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net750 (.A(net750),
    .X(clknet_0_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_0__leaf_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_1__leaf_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net651 (.A(net651),
    .X(clknet_0_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net749 (.A(net749),
    .X(clknet_0_net749));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net749 (.A(clknet_0_net749),
    .X(clknet_1_0__leaf_net749));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net749 (.A(clknet_0_net749),
    .X(clknet_1_1__leaf_net749));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net650 (.A(net650),
    .X(clknet_0_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net650 (.A(clknet_0_net650),
    .X(clknet_1_0__leaf_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net650 (.A(clknet_0_net650),
    .X(clknet_1_1__leaf_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net270 (.A(net270),
    .X(clknet_0_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_0__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net388 (.A(net388),
    .X(clknet_0_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net388 (.A(clknet_0_net388),
    .X(clknet_1_0__leaf_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net388 (.A(clknet_0_net388),
    .X(clknet_1_1__leaf_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net500 (.A(net500),
    .X(clknet_0_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net500 (.A(clknet_0_net500),
    .X(clknet_1_0__leaf_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net500 (.A(clknet_0_net500),
    .X(clknet_1_1__leaf_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net371 (.A(net371),
    .X(clknet_0_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_0__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_1__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net486 (.A(net486),
    .X(clknet_0_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_0__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_1__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net581 (.A(net581),
    .X(clknet_0_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_0__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_1__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net374 (.A(net374),
    .X(clknet_0_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net374 (.A(clknet_0_net374),
    .X(clknet_1_0__leaf_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net374 (.A(clknet_0_net374),
    .X(clknet_1_1__leaf_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net384 (.A(net384),
    .X(clknet_0_net384));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net384 (.A(clknet_0_net384),
    .X(clknet_1_0__leaf_net384));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net384 (.A(clknet_0_net384),
    .X(clknet_1_1__leaf_net384));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net385 (.A(net385),
    .X(clknet_0_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_0__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_1__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net377 (.A(net377),
    .X(clknet_0_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_1__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net373 (.A(net373),
    .X(clknet_0_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net373 (.A(net792),
    .X(clknet_1_1__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net381 (.A(net381),
    .X(clknet_0_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net381 (.A(net788),
    .X(clknet_1_0__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_1__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net507 (.A(net507),
    .X(clknet_0_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_0__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_1__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net513 (.A(net513),
    .X(clknet_0_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_0__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_1__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net491 (.A(net491),
    .X(clknet_0_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_0__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer1 (.A(net752),
    .X(net775));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer2 (.A(net775),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net776),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net775),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(net778),
    .X(net779));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer6 (.A(net787),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net780),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net359),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net782),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net359),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer11 (.A(net88),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net88),
    .X(net786));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer13 (.A(net752),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(clknet_0_net381),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net353),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net789),
    .X(net790));
 sky130_fd_sc_hd__buf_2 rebuffer17 (.A(net790),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(clknet_0_net373),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net451),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net649),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net65),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net67),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net305),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net455),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net320),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net340),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net757),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net485),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net343),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net664),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net453),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net194),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net322),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net527),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net735),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net644),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net286),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net309),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net179),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net342),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net548),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net426),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net647),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net300),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net592),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net180),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net763),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net162),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net545),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net167),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net295),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net280),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net646),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net564),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net740),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net660),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net189),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net62),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net642),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net258),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net169),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net735),
    .X(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_A3 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_Y (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_SCE (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_RESET_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge761_A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_Y (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B_N (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_Y (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge756_A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A4 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_Y (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_SET_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_Y (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_RESET_B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_Y (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_D (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B_N (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge761_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A4 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B_N (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_Y (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B_N (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_Y (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_SCD (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B_N (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_Y (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge761_S0 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A0 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_X (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A0 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_X (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_X (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_Y (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_SCE (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_SCE (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_Y (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_RESET_B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_SCD (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_Y (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A3 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B_N (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_Y (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_D (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B_N (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B1_N (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_SCD (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_DE (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_RESET_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_RESET_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_RESET_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_SCE (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_Y (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_GATE (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_SCD (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B1_N (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_Y (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_D (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_SCD (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_SET_B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_Y (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_D (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SCD (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_SCE (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_SET_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_D (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_SCE (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_SCD (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_SCE (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_SCD (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_X (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_B1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_Y (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A_N (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_B1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_Y (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1_N (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_SCE (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_Y (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_B (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_Q (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SET_B (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_SCE (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_D (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_D (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_Y (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_RESET_B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B1_N (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_X (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge755_SCD (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_SCE (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_Y (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_B_N (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_X (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_X (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_SCE (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_Y (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_DE (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_D (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_RESET_B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_RESET_B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_Y (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B_N (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_B_N (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_Y (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_RESET_B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_Q (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A4 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_SCD (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_X (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_B1_N (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_SCE (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_RESET_B (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_B1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_D (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A3 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B1_N (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_Y (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge756_A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_SCD (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A0 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SCE (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_X (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_Q_N (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SCD (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B_N (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_Q (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_D (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_B1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_Y (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge756_S0 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S0 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_Q_N (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_Q_N (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge755_D (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_B (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_Y (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_B1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_B1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_B_N (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_Y (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SCE (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_DE (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_Y (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_D (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_Y (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_B1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_B (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_X (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_DE (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A4 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_SCD (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_Y (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_SET_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_Q (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_SCE (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_SET_B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_Q_N (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_D (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_Y (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_D (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B1_N (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_Y (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B_N (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_D (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A4 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_B_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_Y (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_RESET_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_Y (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B_N (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A_N (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_Y (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCD (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B_N (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_SET_B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A_N (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_B (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A_N (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_SCE (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A_N (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_B_N (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_B (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_D (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S0 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_S (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_A4 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_N (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A0 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_B1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_B1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_A4 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_A3 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_B1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_B1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_B (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_D (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A_N (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_Q (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B1_N (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_Y (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_SCE (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_Y (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SCE (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_RESET_B (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SCE (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_B1_N (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S0 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1_N (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_Q (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B1_N (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A3 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_RESET_B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_RESET_B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SCD (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SET_B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_X (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SCE (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SET_B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_SET_B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A3 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_SET_B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SCD (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_X (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_Y (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_B1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B_N (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_X (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold57_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B1_N (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_B1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_SET_B (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Y (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_Y (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_B1_N (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A3 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_X (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_S0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_B (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_B (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_B (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_B_N (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_Y (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_SCD (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_RESET_B (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1_N (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_X (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_B1_N (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B1_N (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_Y (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold49_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_Q (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_SCE (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B1_N (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1_N (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_SET_B (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_Y (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap106_A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_Y (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_B1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_B1_N (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B_N (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_SCE (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_Q (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_SET_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SCE (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1_N (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap106_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge761_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_SCD (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A4 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_RESET_B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_SCE (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_SCE (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_S (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B_N (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B1_N (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_B1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_B1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_B1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_B1_N (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B1_N (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCE (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_SCD (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_B1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s762_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s763_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s764_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge758_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s765_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s767_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s766_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s773_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c642_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s772_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s779_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s780_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(clknet_1_0__leaf_net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_SCE (.DIODE(clknet_1_0__leaf_net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(clknet_1_0__leaf_net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net388_X (.DIODE(clknet_1_0__leaf_net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_D (.DIODE(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net377_X (.DIODE(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B_N (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_SET_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_B (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_D (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net688));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net721),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net794),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net794),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net794),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net794),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net794),
    .X(net841));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer25 (.A(net721),
    .X(net843));
 sky130_fd_sc_hd__or2_1 clone26 (.A(net667),
    .B(net715),
    .X(net844));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
