module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net1047;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net1049;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net1053;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net1056;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net1057;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net1058;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire clknet_0_clk;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1048;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1054;
 wire net1055;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net889;
 wire clknet_1_0__leaf_net889;
 wire clknet_1_1__leaf_net889;
 wire clknet_0_net888;
 wire clknet_1_0__leaf_net888;
 wire clknet_1_1__leaf_net888;
 wire clknet_0_net770;
 wire clknet_1_0__leaf_net770;
 wire clknet_1_1__leaf_net770;
 wire clknet_0_net617;
 wire clknet_1_0__leaf_net617;
 wire clknet_1_1__leaf_net617;
 wire clknet_0_net887;
 wire clknet_1_0__leaf_net887;
 wire clknet_1_1__leaf_net887;
 wire clknet_0_net612;
 wire clknet_1_0__leaf_net612;
 wire clknet_1_1__leaf_net612;
 wire clknet_0_net616;
 wire clknet_1_0__leaf_net616;
 wire clknet_1_1__leaf_net616;
 wire clknet_0_net969;
 wire clknet_1_0__leaf_net969;
 wire clknet_1_1__leaf_net969;
 wire clknet_0_net869;
 wire clknet_1_0__leaf_net869;
 wire clknet_1_1__leaf_net869;
 wire clknet_0_net504;
 wire clknet_1_0__leaf_net504;
 wire clknet_1_1__leaf_net504;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net868;
 wire clknet_1_0__leaf_net868;
 wire clknet_1_1__leaf_net868;
 wire clknet_0_net850;
 wire clknet_1_0__leaf_net850;
 wire clknet_1_1__leaf_net850;
 wire clknet_0_net356;
 wire clknet_1_0__leaf_net356;
 wire clknet_1_1__leaf_net356;
 wire clknet_0_net351;
 wire clknet_1_0__leaf_net351;
 wire clknet_1_1__leaf_net351;
 wire clknet_0_net978;
 wire clknet_1_0__leaf_net978;
 wire clknet_1_1__leaf_net978;
 wire clknet_0_net849;
 wire clknet_1_0__leaf_net849;
 wire clknet_1_1__leaf_net849;
 wire clknet_0_net342;
 wire clknet_1_0__leaf_net342;
 wire clknet_1_1__leaf_net342;
 wire clknet_0_net848;
 wire clknet_1_0__leaf_net848;
 wire clknet_1_1__leaf_net848;
 wire clknet_0_net541;
 wire clknet_1_0__leaf_net541;
 wire clknet_1_1__leaf_net541;
 wire clknet_0_net546;
 wire clknet_1_0__leaf_net546;
 wire clknet_1_1__leaf_net546;
 wire clknet_0_net418;
 wire clknet_1_0__leaf_net418;
 wire clknet_1_1__leaf_net418;
 wire clknet_0_net432;
 wire clknet_1_0__leaf_net432;
 wire clknet_1_1__leaf_net432;
 wire clknet_0_net536;
 wire clknet_1_0__leaf_net536;
 wire clknet_1_1__leaf_net536;
 wire clknet_0_net438;
 wire clknet_1_0__leaf_net438;
 wire clknet_1_1__leaf_net438;
 wire clknet_0_net429;
 wire clknet_1_0__leaf_net429;
 wire clknet_1_1__leaf_net429;
 wire clknet_0_net485;
 wire clknet_1_0__leaf_net485;
 wire clknet_1_1__leaf_net485;
 wire clknet_0_net464;
 wire clknet_1_0__leaf_net464;
 wire clknet_1_1__leaf_net464;
 wire clknet_0_net427;
 wire clknet_1_0__leaf_net427;
 wire clknet_1_1__leaf_net427;
 wire clknet_0_net445;
 wire clknet_1_0__leaf_net445;
 wire clknet_1_1__leaf_net445;
 wire clknet_0_net967;
 wire clknet_1_0__leaf_net967;
 wire clknet_1_1__leaf_net967;
 wire clknet_0_net503;
 wire clknet_1_0__leaf_net503;
 wire clknet_1_1__leaf_net503;
 wire clknet_0_net425;
 wire clknet_1_0__leaf_net425;
 wire clknet_1_1__leaf_net425;
 wire clknet_0_net430;
 wire clknet_1_0__leaf_net430;
 wire clknet_1_1__leaf_net430;
 wire clknet_0_net417;
 wire clknet_1_0__leaf_net417;
 wire clknet_1_1__leaf_net417;
 wire clknet_0_net1002;
 wire clknet_1_0__leaf_net1002;
 wire clknet_1_1__leaf_net1002;
 wire clknet_0_net190;
 wire clknet_1_0__leaf_net190;
 wire clknet_1_1__leaf_net190;
 wire clknet_0_net993;
 wire clknet_1_0__leaf_net993;
 wire clknet_1_1__leaf_net993;
 wire clknet_0_net992;
 wire clknet_1_0__leaf_net992;
 wire clknet_1_1__leaf_net992;
 wire clknet_0_net832;
 wire clknet_1_0__leaf_net832;
 wire clknet_1_1__leaf_net832;
 wire clknet_0_net371;
 wire clknet_1_0__leaf_net371;
 wire clknet_1_1__leaf_net371;
 wire clknet_0_net374;
 wire clknet_1_0__leaf_net374;
 wire clknet_1_1__leaf_net374;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net986;
 wire clknet_1_0__leaf_net986;
 wire clknet_1_1__leaf_net986;
 wire clknet_0_net36;
 wire clknet_1_0__leaf_net36;
 wire clknet_1_1__leaf_net36;
 wire clknet_0_net38;
 wire clknet_1_0__leaf_net38;
 wire clknet_1_1__leaf_net38;
 wire clknet_0_net35;
 wire clknet_1_0__leaf_net35;
 wire clknet_1_1__leaf_net35;
 wire clknet_0_net39;
 wire clknet_1_0__leaf_net39;
 wire clknet_1_1__leaf_net39;
 wire clknet_0_net998;
 wire clknet_1_0__leaf_net998;
 wire clknet_1_1__leaf_net998;
 wire clknet_0_net304;
 wire clknet_1_0__leaf_net304;
 wire clknet_1_1__leaf_net304;
 wire clknet_0_net516;
 wire clknet_1_0__leaf_net516;
 wire clknet_1_1__leaf_net516;
 wire clknet_0_net172;
 wire clknet_1_0__leaf_net172;
 wire clknet_1_1__leaf_net172;
 wire clknet_0_net175;
 wire clknet_1_0__leaf_net175;
 wire clknet_1_1__leaf_net175;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net176;
 wire clknet_1_0__leaf_net176;
 wire clknet_1_1__leaf_net176;
 wire clknet_0_net168;
 wire clknet_1_0__leaf_net168;
 wire clknet_1_1__leaf_net168;
 wire clknet_0_net961;
 wire clknet_1_0__leaf_net961;
 wire clknet_1_1__leaf_net961;
 wire clknet_0_net167;
 wire clknet_1_0__leaf_net167;
 wire clknet_1_1__leaf_net167;
 wire clknet_0_net24;
 wire clknet_1_0__leaf_net24;
 wire clknet_1_1__leaf_net24;
 wire clknet_0_net25;
 wire clknet_1_0__leaf_net25;
 wire clknet_1_1__leaf_net25;
 wire clknet_0_net54;
 wire clknet_1_0__leaf_net54;
 wire clknet_1_1__leaf_net54;
 wire clknet_0_net19;
 wire clknet_1_0__leaf_net19;
 wire clknet_1_1__leaf_net19;
 wire clknet_0_net1010;
 wire clknet_1_0__leaf_net1010;
 wire clknet_1_1__leaf_net1010;
 wire clknet_0_net22;
 wire clknet_1_0__leaf_net22;
 wire clknet_1_1__leaf_net22;
 wire clknet_0_net140;
 wire clknet_1_0__leaf_net140;
 wire clknet_1_1__leaf_net140;
 wire clknet_0_net29;
 wire clknet_1_0__leaf_net29;
 wire clknet_1_1__leaf_net29;
 wire clknet_0_net34;
 wire clknet_1_0__leaf_net34;
 wire clknet_1_1__leaf_net34;
 wire clknet_0_net30;
 wire clknet_1_0__leaf_net30;
 wire clknet_1_1__leaf_net30;
 wire clknet_0_net769;
 wire clknet_1_0__leaf_net769;
 wire clknet_1_1__leaf_net769;
 wire clknet_0_net12;
 wire clknet_1_0__leaf_net12;
 wire clknet_1_1__leaf_net12;
 wire clknet_0_net16;
 wire clknet_1_0__leaf_net16;
 wire clknet_1_1__leaf_net16;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net303;
 wire clknet_1_0__leaf_net303;
 wire clknet_1_1__leaf_net303;
 wire clknet_0_net169;
 wire clknet_1_0__leaf_net169;
 wire clknet_1_1__leaf_net169;
 wire clknet_0_net157;
 wire clknet_1_0__leaf_net157;
 wire clknet_1_1__leaf_net157;
 wire clknet_0_net1008;
 wire clknet_1_0__leaf_net1008;
 wire clknet_1_1__leaf_net1008;
 wire clknet_0_net130;
 wire clknet_1_0__leaf_net130;
 wire clknet_1_1__leaf_net130;
 wire clknet_0_net111;
 wire clknet_1_0__leaf_net111;
 wire clknet_1_1__leaf_net111;
 wire clknet_0_net110;
 wire clknet_1_0__leaf_net110;
 wire clknet_1_1__leaf_net110;
 wire net17;
 wire net23;
 wire net133;
 wire net152;
 wire net450;
 wire net570;
 wire net962;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;

 sky130_fd_sc_hd__nand2_1 c100 (.A(net20),
    .B(net27),
    .Y(net37));
 sky130_fd_sc_hd__mux4_4 c101 (.A0(clknet_1_1__leaf_net35),
    .A1(clknet_1_0__leaf_net36),
    .A2(net37),
    .A3(net28),
    .S0(net927),
    .S1(net33),
    .X(net38));
 sky130_fd_sc_hd__o211a_4 c102 (.A1(net37),
    .A2(net928),
    .B1(net33),
    .C1(clknet_1_0__leaf_net35),
    .X(net39));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net26),
    .A1(clknet_1_1__leaf_net36),
    .A2(net33),
    .A3(net1014),
    .S0(clknet_1_0__leaf_net39),
    .S1(clknet_1_1__leaf_net34),
    .X(net40));
 sky130_fd_sc_hd__sdfrbp_2 c104 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_0__leaf_net39),
    .RESET_B(clknet_1_1__leaf_net34),
    .SCD(net33),
    .SCE(clknet_1_1__leaf_net25),
    .Q(net42),
    .Q_N(net41));
 sky130_fd_sc_hd__inv_4 c105 (.A(net816),
    .Y(net43));
 sky130_fd_sc_hd__o211ai_2 c106 (.A1(net947),
    .A2(clknet_1_1__leaf_net39),
    .B1(net31),
    .C1(net827),
    .Y(net44));
 sky130_fd_sc_hd__sdfrbp_2 c107 (.CLK(clknet_4_13_0_clk),
    .D(net31),
    .RESET_B(net1075),
    .SCD(net1014),
    .SCE(net725),
    .Q(net997),
    .Q_N(net45));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(clknet_1_0__leaf_net35),
    .A1(net1052),
    .A2(clknet_1_0__leaf_net30),
    .A3(net33),
    .S0(net28),
    .X(net46));
 sky130_fd_sc_hd__sdfbbn_2 c109 (.CLK_N(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net39),
    .RESET_B(net997),
    .SCD(net32),
    .SCE(net41),
    .SET_B(net725),
    .Q(net48),
    .Q_N(net47));
 sky130_fd_sc_hd__clkbuf_1 c110 (.A(net654),
    .X(net49));
 sky130_fd_sc_hd__nand2_2 c111 (.A(net920),
    .B(clknet_1_0__leaf_net24),
    .Y(net50));
 sky130_fd_sc_hd__and3b_1 c112 (.A_N(net9),
    .B(net11),
    .C(net45),
    .X(net51));
 sky130_fd_sc_hd__and2b_1 c113 (.A_N(net43),
    .B(net920),
    .X(net52));
 sky130_fd_sc_hd__or2_1 c114 (.A(net926),
    .B(net45),
    .X(net53));
 sky130_fd_sc_hd__and2_1 c115 (.A(clknet_1_1__leaf_net24),
    .B(net43),
    .X(net54));
 sky130_fd_sc_hd__nand2b_2 c116 (.A_N(net51),
    .B(net52),
    .Y(net55));
 sky130_fd_sc_hd__nand2b_1 c117 (.A_N(net917),
    .B(net43),
    .Y(net56));
 sky130_fd_sc_hd__o211a_1 c118 (.A1(net49),
    .A2(net55),
    .B1(net52),
    .C1(net1014),
    .X(net57));
 sky130_fd_sc_hd__sdfrtn_1 c119 (.CLK_N(clknet_4_15_0_clk),
    .D(net53),
    .RESET_B(net1070),
    .SCD(net926),
    .SCE(net55),
    .Q(net58));
 sky130_fd_sc_hd__nor2b_1 c120 (.A(net32),
    .B_N(net1042),
    .Y(net59));
 sky130_fd_sc_hd__nor3_1 c121 (.A(net59),
    .B(net1045),
    .C(net1042),
    .Y(net60));
 sky130_fd_sc_hd__sdfrtp_1 c122 (.CLK(clknet_4_15_0_clk),
    .D(net52),
    .RESET_B(clknet_1_0__leaf_net54),
    .SCD(net60),
    .SCE(net55),
    .Q(net61));
 sky130_fd_sc_hd__inv_6 c123 (.A(net654),
    .Y(net974));
 sky130_fd_sc_hd__nand2_1 c124 (.A(net3),
    .B(net51),
    .Y(net62));
 sky130_fd_sc_hd__o221ai_1 c125 (.A1(net62),
    .A2(net59),
    .B1(net1042),
    .B2(net1014),
    .C1(net1085),
    .Y(net63));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net61),
    .A1(net902),
    .A2(net921),
    .A3(net1042),
    .S0(net1044),
    .S1(net11),
    .X(net64));
 sky130_fd_sc_hd__o221a_1 c127 (.A1(net56),
    .A2(net59),
    .B1(net1042),
    .B2(net902),
    .C1(net61),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(clknet_1_0__leaf_net38),
    .A1(net1042),
    .A2(net65),
    .A3(net810),
    .S0(net813),
    .S1(net827),
    .X(net66));
 sky130_fd_sc_hd__inv_1 c129 (.A(net816),
    .Y(net67));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net50),
    .A1(net67),
    .A2(net62),
    .A3(net65),
    .S0(net51),
    .S1(net1042),
    .X(net68));
 sky130_fd_sc_hd__sdfbbn_1 c131 (.CLK_N(clknet_4_15_0_clk),
    .D(net62),
    .RESET_B(net1042),
    .SCD(clknet_1_1__leaf_net54),
    .SCE(net810),
    .SET_B(net828),
    .Q(net70),
    .Q_N(net69));
 sky130_fd_sc_hd__and2_2 c132 (.A(net932),
    .B(net957),
    .X(net71));
 sky130_fd_sc_hd__nand3b_4 c133 (.A_N(net907),
    .B(net954),
    .C(net905),
    .Y(net72));
 sky130_fd_sc_hd__nand2b_2 c134 (.A_N(net1041),
    .B(net907),
    .Y(net73));
 sky130_fd_sc_hd__o211ai_2 c135 (.A1(net932),
    .A2(net908),
    .B1(net1041),
    .C1(net921),
    .Y(net74));
 sky130_fd_sc_hd__or3_2 c136 (.A(net909),
    .B(net958),
    .C(net1041),
    .X(net75));
 sky130_fd_sc_hd__or3b_2 c137 (.A(net75),
    .B(net899),
    .C_N(net902),
    .X(net76));
 sky130_fd_sc_hd__and2_1 c138 (.A(net903),
    .B(net900),
    .X(net77));
 sky130_fd_sc_hd__inv_12 c139 (.A(net765),
    .Y(net78));
 sky130_fd_sc_hd__nor2_1 c140 (.A(net954),
    .B(net910),
    .Y(net79));
 sky130_fd_sc_hd__o221ai_4 c141 (.A1(net75),
    .A2(net73),
    .B1(net908),
    .B2(net957),
    .C1(net959),
    .Y(net80));
 sky130_fd_sc_hd__or3_4 c142 (.A(net958),
    .B(net1043),
    .C(net1041),
    .X(net81));
 sky130_fd_sc_hd__inv_4 c143 (.A(net765),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 c144 (.A(net749),
    .Y(net83));
 sky130_fd_sc_hd__mux4_1 c145 (.A0(net901),
    .A1(net1040),
    .A2(net83),
    .A3(net73),
    .S0(net80),
    .S1(net959),
    .X(net84));
 sky130_fd_sc_hd__or2_2 c146 (.A(net1040),
    .B(net763),
    .X(net85));
 sky130_fd_sc_hd__or2_4 c147 (.A(net82),
    .B(net905),
    .X(net86));
 sky130_fd_sc_hd__or3_1 c148 (.A(net83),
    .B(net85),
    .C(net86),
    .X(net87));
 sky130_fd_sc_hd__inv_4 c149 (.A(net765),
    .Y(net88));
 sky130_fd_sc_hd__nand3b_1 c150 (.A_N(net905),
    .B(net78),
    .C(net83),
    .Y(net89));
 sky130_fd_sc_hd__nand3_1 c151 (.A(net74),
    .B(net1083),
    .C(net86),
    .Y(net90));
 sky130_fd_sc_hd__o211a_1 c152 (.A1(net88),
    .A2(net78),
    .B1(net79),
    .C1(net83),
    .X(net91));
 sky130_fd_sc_hd__sdfrtp_4 c153 (.CLK(clknet_4_5_0_clk),
    .D(net91),
    .RESET_B(net90),
    .SCD(net86),
    .SCE(net81),
    .Q(net92));
 sky130_fd_sc_hd__or2_1 c154 (.A(net936),
    .B(net900),
    .X(net93));
 sky130_fd_sc_hd__or2_1 c155 (.A(net910),
    .B(net914),
    .X(net94));
 sky130_fd_sc_hd__nor3b_2 c156 (.A(net922),
    .B(net83),
    .C_N(net1034),
    .Y(net95));
 sky130_fd_sc_hd__nand3b_4 c157 (.A_N(net911),
    .B(net922),
    .C(net1034),
    .Y(net96));
 sky130_fd_sc_hd__and2b_1 c158 (.A_N(net93),
    .B(net1034),
    .X(net97));
 sky130_fd_sc_hd__nor3_1 c159 (.A(net93),
    .B(net933),
    .C(net1034),
    .Y(net98));
 sky130_fd_sc_hd__o211ai_1 c160 (.A1(net97),
    .A2(net1031),
    .B1(net927),
    .C1(net1034),
    .Y(net99));
 sky130_fd_sc_hd__o211a_1 c161 (.A1(net908),
    .A2(net935),
    .B1(net1031),
    .C1(net1034),
    .X(net100));
 sky130_fd_sc_hd__inv_6 c162 (.A(net759),
    .Y(net101));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net959),
    .A1(net908),
    .A2(net101),
    .A3(net92),
    .S0(net1031),
    .S1(net1034),
    .X(net102));
 sky130_fd_sc_hd__o211a_1 c164 (.A1(net97),
    .A2(net899),
    .B1(net1031),
    .C1(net1035),
    .X(net103));
 sky130_fd_sc_hd__o211ai_1 c165 (.A1(net916),
    .A2(net103),
    .B1(net99),
    .C1(net1034),
    .Y(net104));
 sky130_fd_sc_hd__clkbuf_1 c166 (.A(net759),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 c167 (.A(net771),
    .X(net106));
 sky130_fd_sc_hd__sdfbbp_1 c168 (.CLK(clknet_4_7_0_clk),
    .D(net105),
    .RESET_B(net100),
    .SCD(net101),
    .SCE(net78),
    .SET_B(net1035),
    .Q(net108),
    .Q_N(net107));
 sky130_fd_sc_hd__nand3_2 c169 (.A(net925),
    .B(net1034),
    .C(net765),
    .Y(net109));
 sky130_fd_sc_hd__o221a_2 c170 (.A1(net106),
    .A2(net101),
    .B1(net98),
    .B2(net1035),
    .C1(net765),
    .X(net110));
 sky130_fd_sc_hd__o221a_1 c171 (.A1(net106),
    .A2(net109),
    .B1(net107),
    .B2(net96),
    .C1(net1035),
    .X(net111));
 sky130_fd_sc_hd__sdfbbn_1 c172 (.CLK_N(clknet_4_7_0_clk),
    .D(net96),
    .RESET_B(net105),
    .SCD(clknet_1_0__leaf_net110),
    .SCE(net109),
    .SET_B(net1035),
    .Q(net113),
    .Q_N(net112));
 sky130_fd_sc_hd__sdfbbn_1 c173 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net110),
    .RESET_B(net108),
    .SCD(net1096),
    .SCE(net1035),
    .SET_B(net106),
    .Q(net115),
    .Q_N(net114));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(clknet_1_0__leaf_net111),
    .A1(net105),
    .A2(net101),
    .A3(net106),
    .S0(net112),
    .S1(net763),
    .X(net116));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net99),
    .A1(clknet_1_0__leaf_net110),
    .A2(net922),
    .A3(net112),
    .S0(net109),
    .S1(net829),
    .X(net117));
 sky130_fd_sc_hd__inv_2 c176 (.A(net759),
    .Y(net118));
 sky130_fd_sc_hd__or2_2 c177 (.A(net108),
    .B(net114),
    .X(net119));
 sky130_fd_sc_hd__nor2_1 c178 (.A(net119),
    .B(net113),
    .Y(net120));
 sky130_fd_sc_hd__nor2b_1 c179 (.A(net942),
    .B_N(net0),
    .Y(net121));
 sky130_fd_sc_hd__and2b_1 c180 (.A_N(net956),
    .B(net952),
    .X(net122));
 sky130_fd_sc_hd__nand2b_1 c181 (.A_N(net83),
    .B(net122),
    .Y(net123));
 sky130_fd_sc_hd__nor3_2 c182 (.A(net938),
    .B(net123),
    .C(net119),
    .Y(net124));
 sky130_fd_sc_hd__buf_4 c183 (.A(net745),
    .X(net125));
 sky130_fd_sc_hd__or2_4 c184 (.A(net109),
    .B(net125),
    .X(net1000));
 sky130_fd_sc_hd__inv_1 c185 (.A(net820),
    .Y(net126));
 sky130_fd_sc_hd__clkbuf_4 c186 (.A(net820),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 c187 (.A(net763),
    .X(net128));
 sky130_fd_sc_hd__nor2b_1 c188 (.A(net126),
    .B_N(net123),
    .Y(net129));
 sky130_fd_sc_hd__mux4_4 c189 (.A0(net120),
    .A1(net106),
    .A2(net952),
    .A3(net128),
    .S0(net107),
    .S1(net127),
    .X(net130));
 sky130_fd_sc_hd__and3b_1 c190 (.A_N(net128),
    .B(net127),
    .C(net1039),
    .X(net131));
 sky130_fd_sc_hd__and2_1 c191 (.A(net131),
    .B(net127),
    .X(net132));
 sky130_fd_sc_hd__clkinv_2 c214_2 (.A(net771),
    .Y(net1047));
 sky130_fd_sc_hd__mux4_4 c193 (.A0(net125),
    .A1(net77),
    .A2(net124),
    .A3(net132),
    .S0(net914),
    .S1(net112),
    .X(net134));
 sky130_fd_sc_hd__inv_4 c194 (.A(net763),
    .Y(net135));
 sky130_fd_sc_hd__or2_2 c195 (.A(net126),
    .B(net830),
    .X(net136));
 sky130_fd_sc_hd__mux4_2 c196 (.A0(net1046),
    .A1(net944),
    .A2(net136),
    .A3(net83),
    .S0(net1031),
    .S1(net1000),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net132),
    .A1(net122),
    .A2(net136),
    .A3(net127),
    .S0(net135),
    .S1(net830),
    .X(net138));
 sky130_fd_sc_hd__and3b_1 c198 (.A_N(net92),
    .B(net115),
    .C(net1039),
    .X(net139));
 sky130_fd_sc_hd__o221ai_2 c199 (.A1(net139),
    .A2(clknet_1_0__leaf_net22),
    .B1(net1041),
    .B2(net136),
    .C1(net96),
    .Y(net140));
 sky130_fd_sc_hd__buf_6 c200 (.A(net721),
    .X(net141));
 sky130_fd_sc_hd__buf_6 c201 (.A(net810),
    .X(net142));
 sky130_fd_sc_hd__inv_6 c202 (.A(net789),
    .Y(net996));
 sky130_fd_sc_hd__and2_2 c203 (.A(net141),
    .B(net740),
    .X(net143));
 sky130_fd_sc_hd__inv_1 c204 (.A(net790),
    .Y(net144));
 sky130_fd_sc_hd__and2b_1 c205 (.A_N(net918),
    .B(net136),
    .X(net145));
 sky130_fd_sc_hd__nand3b_4 c206 (.A_N(net145),
    .B(net127),
    .C(net143),
    .Y(net146));
 sky130_fd_sc_hd__clkinv_4 c207 (.A(net777),
    .Y(net147));
 sky130_fd_sc_hd__nand3_4 c208 (.A(net949),
    .B(net147),
    .C(net830),
    .Y(net1003));
 sky130_fd_sc_hd__clkbuf_2 c209 (.A(net721),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 c210 (.A(net743),
    .X(net149));
 sky130_fd_sc_hd__nand3b_4 c211 (.A_N(net136),
    .B(net145),
    .C(net148),
    .Y(net988));
 sky130_fd_sc_hd__sdfrtp_2 c212 (.CLK(clknet_4_12_0_clk),
    .D(net147),
    .RESET_B(net141),
    .SCD(net146),
    .SCE(net1022),
    .Q(net150));
 sky130_fd_sc_hd__o211a_1 c213 (.A1(net1003),
    .A2(net115),
    .B1(net144),
    .C1(net830),
    .X(net151));
 sky130_fd_sc_hd__clkinv_8 c79_4 (.A(net771),
    .Y(net1049));
 sky130_fd_sc_hd__inv_8 c215 (.A(net788),
    .Y(net153));
 sky130_fd_sc_hd__o211a_2 c216 (.A1(net148),
    .A2(net150),
    .B1(net149),
    .C1(net151),
    .X(net1004));
 sky130_fd_sc_hd__o211a_1 c217 (.A1(net150),
    .A2(net146),
    .B1(net919),
    .C1(net1086),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net1048),
    .A1(net149),
    .A2(net146),
    .A3(net141),
    .S0(net153),
    .S1(net721),
    .X(net155));
 sky130_fd_sc_hd__mux4_2 c219 (.A0(net988),
    .A1(net1004),
    .A2(net136),
    .A3(net146),
    .S0(net721),
    .S1(clknet_1_1__leaf_net832),
    .X(net156));
 sky130_fd_sc_hd__nand3_4 c220 (.A(net903),
    .B(net127),
    .C(clknet_1_1__leaf_net12),
    .Y(net157));
 sky130_fd_sc_hd__nor2b_2 c221 (.A(clknet_1_1__leaf_net29),
    .B_N(net917),
    .Y(net1008));
 sky130_fd_sc_hd__o211a_4 c222 (.A1(net902),
    .A2(net28),
    .B1(clknet_1_1__leaf_net157),
    .C1(net988),
    .X(net158));
 sky130_fd_sc_hd__buf_2 c223 (.A(net813),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd1_1 c224 (.A(net804),
    .X(net160));
 sky130_fd_sc_hd__inv_1 c225 (.A(net760),
    .Y(net161));
 sky130_fd_sc_hd__or2b_2 c226 (.A(clknet_1_1__leaf_net12),
    .B_N(net1039),
    .X(net162));
 sky130_fd_sc_hd__sdfsbp_1 c227 (.CLK(clknet_4_15_0_clk),
    .D(clknet_1_1__leaf_net25),
    .SCD(net926),
    .SCE(clknet_1_1__leaf_net162),
    .SET_B(clknet_1_0__leaf_net160),
    .Q(net164),
    .Q_N(net163));
 sky130_fd_sc_hd__o211ai_4 c228 (.A1(clknet_1_0__leaf_net30),
    .A2(net1003),
    .B1(clknet_1_0__leaf_net25),
    .C1(net14),
    .Y(net165));
 sky130_fd_sc_hd__o211ai_1 c229 (.A1(net917),
    .A2(clknet_1_0__leaf_net29),
    .B1(net163),
    .C1(net2),
    .Y(net166));
 sky130_fd_sc_hd__o221ai_4 c230 (.A1(net143),
    .A2(clknet_1_1__leaf_net19),
    .B1(net997),
    .B2(clknet_1_0__leaf_net160),
    .C1(net28),
    .Y(net167));
 sky130_fd_sc_hd__o221ai_2 c231 (.A1(net28),
    .A2(clknet_1_0__leaf_net160),
    .B1(net47),
    .B2(clknet_1_1__leaf_net12),
    .C1(net1003),
    .Y(net168));
 sky130_fd_sc_hd__nand2b_2 c232 (.A_N(clknet_1_1__leaf_net162),
    .B(clknet_1_1__leaf_net769),
    .Y(net169));
 sky130_fd_sc_hd__sdfsbp_2 c233 (.CLK(clknet_4_15_0_clk),
    .D(clknet_1_0__leaf_net1008),
    .SCD(net127),
    .SCE(clknet_1_0__leaf_net167),
    .SET_B(clknet_1_1__leaf_net769),
    .Q(net171),
    .Q_N(net170));
 sky130_fd_sc_hd__buf_2 c234 (.A(net804),
    .X(net172));
 sky130_fd_sc_hd__sdfbbp_1 c235 (.CLK(clknet_4_12_0_clk),
    .D(net917),
    .RESET_B(clknet_1_0__leaf_net157),
    .SCD(net1014),
    .SCE(net948),
    .SET_B(net1065),
    .Q(net174),
    .Q_N(net173));
 sky130_fd_sc_hd__mux4_2 c236 (.A0(clknet_1_0__leaf_net157),
    .A1(clknet_1_1__leaf_net22),
    .A2(net171),
    .A3(clknet_1_1__leaf_net162),
    .S0(net1044),
    .S1(clknet_1_0__leaf_net172),
    .X(net175));
 sky130_fd_sc_hd__o221ai_2 c237 (.A1(net953),
    .A2(net161),
    .B1(clknet_1_1__leaf_net160),
    .B2(net173),
    .C1(net170),
    .Y(net176));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net1055),
    .A1(net174),
    .A2(clknet_1_1__leaf_net167),
    .A3(clknet_1_1__leaf_net160),
    .S0(clknet_1_1__leaf_net169),
    .S1(clknet_1_0__leaf_net176),
    .X(net177));
 sky130_fd_sc_hd__sdfstp_1 c239 (.CLK(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net172),
    .SCD(net164),
    .SCE(clknet_1_1__leaf_net167),
    .SET_B(net1071),
    .Q(net178));
 sky130_fd_sc_hd__nand2_1 c240 (.A(net174),
    .B(net171),
    .Y(net179));
 sky130_fd_sc_hd__o221a_1 c241 (.A1(net179),
    .A2(net178),
    .B1(net159),
    .B2(net1044),
    .C1(net779),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_2 c242 (.A(net798),
    .X(net180));
 sky130_fd_sc_hd__or3b_1 c243 (.A(net64),
    .B(net997),
    .C_N(net983),
    .X(net181));
 sky130_fd_sc_hd__and2_1 c244 (.A(clknet_1_1__leaf_net176),
    .B(clknet_1_0__leaf_net168),
    .X(net182));
 sky130_fd_sc_hd__and3_1 c245 (.A(net14),
    .B(net70),
    .C(net64),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd1_1 c246 (.A(net798),
    .X(net1001));
 sky130_fd_sc_hd__nor3b_2 c247 (.A(clknet_1_1__leaf_net160),
    .B(net48),
    .C_N(net1001),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 c248 (.A(net793),
    .Y(net185));
 sky130_fd_sc_hd__mux4_2 c249 (.A0(net164),
    .A1(clknet_1_0__leaf_net54),
    .A2(net180),
    .A3(net912),
    .S0(clknet_1_0__leaf_net160),
    .S1(net14),
    .X(net186));
 sky130_fd_sc_hd__clkinv_8 c250 (.A(net789),
    .Y(net187));
 sky130_fd_sc_hd__mux4_4 c251 (.A0(net153),
    .A1(net187),
    .A2(net163),
    .A3(net1042),
    .S0(clknet_1_1__leaf_net54),
    .S1(net185),
    .X(net188));
 sky130_fd_sc_hd__o211a_1 c252 (.A1(clknet_1_1__leaf_net54),
    .A2(net69),
    .B1(net187),
    .C1(clknet_1_0__leaf_net1002),
    .X(net189));
 sky130_fd_sc_hd__and3b_2 c253 (.A_N(net187),
    .B(net1038),
    .C(clknet_1_0__leaf_net1002),
    .X(net190));
 sky130_fd_sc_hd__dfbbn_1 c254 (.CLK_N(clknet_4_14_0_clk),
    .D(net1079),
    .RESET_B(net185),
    .SET_B(net183),
    .Q(net192),
    .Q_N(net191));
 sky130_fd_sc_hd__or3_4 c255 (.A(net14),
    .B(net974),
    .C(net787),
    .X(net970));
 sky130_fd_sc_hd__o221ai_2 c256 (.A1(net184),
    .A2(clknet_1_0__leaf_net190),
    .B1(net187),
    .B2(net970),
    .C1(clknet_1_0__leaf_net1002),
    .Y(net193));
 sky130_fd_sc_hd__mux4_4 c257 (.A0(clknet_1_1__leaf_net190),
    .A1(net64),
    .A2(net970),
    .A3(net47),
    .S0(net183),
    .S1(clknet_1_1__leaf_net1002),
    .X(net194));
 sky130_fd_sc_hd__and3b_1 c258 (.A_N(net70),
    .B(net77),
    .C(net787),
    .X(net195));
 sky130_fd_sc_hd__buf_4 c259 (.A(net805),
    .X(net998));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net195),
    .A1(net192),
    .A2(net970),
    .A3(net187),
    .S0(net47),
    .S1(net18),
    .X(net196));
 sky130_fd_sc_hd__mux4_2 c261 (.A0(net923),
    .A1(net195),
    .A2(net970),
    .A3(net187),
    .S0(net805),
    .S1(clknet_1_1__leaf_net1002),
    .X(net197));
 sky130_fd_sc_hd__mux4_2 c262 (.A0(net191),
    .A1(clknet_1_0__leaf_net190),
    .A2(clknet_1_0__leaf_net998),
    .A3(net187),
    .S0(net999),
    .S1(net805),
    .X(net993));
 sky130_fd_sc_hd__o221a_4 c263 (.A1(net181),
    .A2(clknet_1_1__leaf_net190),
    .B1(net48),
    .B2(net970),
    .C1(clknet_1_0__leaf_net993),
    .X(net198));
 sky130_fd_sc_hd__nand2b_4 c264 (.A_N(net899),
    .B(net957),
    .Y(net199));
 sky130_fd_sc_hd__and2_4 c265 (.A(net958),
    .B(net85),
    .X(net200));
 sky130_fd_sc_hd__buf_6 c266 (.A(net735),
    .X(net201));
 sky130_fd_sc_hd__nand2b_1 c267 (.A_N(net905),
    .B(net79),
    .Y(net202));
 sky130_fd_sc_hd__and2_1 c268 (.A(net202),
    .B(net201),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 c269 (.A(net765),
    .X(net204));
 sky130_fd_sc_hd__inv_6 c270 (.A(net748),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 c271 (.A(net735),
    .Y(net206));
 sky130_fd_sc_hd__inv_12 c272 (.A(net749),
    .Y(net207));
 sky130_fd_sc_hd__buf_1 c273 (.A(net962),
    .X(net208));
 sky130_fd_sc_hd__or3b_1 c274 (.A(net202),
    .B(net207),
    .C_N(net943),
    .X(net209));
 sky130_fd_sc_hd__inv_6 c275 (.A(net751),
    .Y(net210));
 sky130_fd_sc_hd__nor3b_1 c276 (.A(net89),
    .B(net208),
    .C_N(net207),
    .Y(net211));
 sky130_fd_sc_hd__buf_2 c277 (.A(net775),
    .X(net212));
 sky130_fd_sc_hd__clkinv_4 c278 (.A(net751),
    .Y(net213));
 sky130_fd_sc_hd__inv_4 c279 (.A(net734),
    .Y(net214));
 sky130_fd_sc_hd__and3_4 c280 (.A(net199),
    .B(net207),
    .C(net213),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c281 (.A0(net214),
    .A1(net212),
    .A2(net210),
    .A3(net907),
    .S0(net213),
    .S1(net207),
    .X(net216));
 sky130_fd_sc_hd__sdfbbn_2 c282 (.CLK_N(clknet_4_5_0_clk),
    .D(net209),
    .RESET_B(net216),
    .SCD(net215),
    .SCE(net213),
    .SET_B(net212),
    .Q(net218),
    .Q_N(net217));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net904),
    .A1(net213),
    .A2(net215),
    .A3(net217),
    .S0(net200),
    .S1(net209),
    .X(net219));
 sky130_fd_sc_hd__sdfbbn_2 c284 (.CLK_N(clknet_4_5_0_clk),
    .D(net202),
    .RESET_B(net214),
    .SCD(net217),
    .SCE(net200),
    .SET_B(net1073),
    .Q(net221),
    .Q_N(net220));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net221),
    .A1(net87),
    .A2(net199),
    .A3(net212),
    .S0(net215),
    .S1(net834),
    .X(net222));
 sky130_fd_sc_hd__nand2b_1 c286 (.A_N(net95),
    .B(net215),
    .Y(net223));
 sky130_fd_sc_hd__nor2b_4 c287 (.A(net929),
    .B_N(net914),
    .Y(net224));
 sky130_fd_sc_hd__mux4_1 c288 (.A0(net224),
    .A1(net79),
    .A2(net98),
    .A3(net100),
    .S0(net1034),
    .S1(net765),
    .X(net225));
 sky130_fd_sc_hd__buf_1 c289 (.A(net768),
    .X(net226));
 sky130_fd_sc_hd__or2b_1 c290 (.A(net79),
    .B_N(net829),
    .X(net227));
 sky130_fd_sc_hd__nand2_1 c291 (.A(net93),
    .B(net86),
    .Y(net228));
 sky130_fd_sc_hd__or2b_2 c292 (.A(net226),
    .B_N(net224),
    .X(net229));
 sky130_fd_sc_hd__or3b_2 c293 (.A(net933),
    .B(net212),
    .C_N(net1036),
    .X(net230));
 sky130_fd_sc_hd__and2b_1 c294 (.A_N(net101),
    .B(net933),
    .X(net231));
 sky130_fd_sc_hd__nand2b_1 c295 (.A_N(net231),
    .B(net212),
    .Y(net232));
 sky130_fd_sc_hd__or2b_2 c296 (.A(net231),
    .B_N(net229),
    .X(net233));
 sky130_fd_sc_hd__o211ai_4 c297 (.A1(net232),
    .A2(net230),
    .B1(net915),
    .C1(net1036),
    .Y(net1006));
 sky130_fd_sc_hd__o221a_2 c298 (.A1(net227),
    .A2(net927),
    .B1(net229),
    .B2(net224),
    .C1(net1036),
    .X(net234));
 sky130_fd_sc_hd__inv_4 c299 (.A(net1090),
    .Y(net235));
 sky130_fd_sc_hd__clkinv_4 c300 (.A(net768),
    .Y(net236));
 sky130_fd_sc_hd__o221a_4 c301 (.A1(net235),
    .A2(net229),
    .B1(net92),
    .B2(net236),
    .C1(net1036),
    .X(net237));
 sky130_fd_sc_hd__buf_1 c302 (.A(net775),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 c303 (.A(net734),
    .X(net239));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net100),
    .A1(net236),
    .A2(net233),
    .A3(net217),
    .S0(net231),
    .S1(net224),
    .X(net240));
 sky130_fd_sc_hd__and2_1 c305 (.A(net218),
    .B(net812),
    .X(net241));
 sky130_fd_sc_hd__or3b_1 c306 (.A(net241),
    .B(net1036),
    .C_N(net812),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net242),
    .A1(net237),
    .A2(net238),
    .A3(net235),
    .S0(net1019),
    .S1(net224),
    .X(net243));
 sky130_fd_sc_hd__nand3_2 c308 (.A(net939),
    .B(net224),
    .C(net1041),
    .Y(net244));
 sky130_fd_sc_hd__or3_1 c309 (.A(net235),
    .B(net118),
    .C(net831),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 c310 (.A(net768),
    .X(net246));
 sky130_fd_sc_hd__inv_4 c311 (.A(net748),
    .Y(net247));
 sky130_fd_sc_hd__buf_1 c312 (.A(net768),
    .X(net248));
 sky130_fd_sc_hd__mux4_4 c313 (.A0(net248),
    .A1(net247),
    .A2(clknet_1_0__leaf_net111),
    .A3(net224),
    .S0(net1019),
    .S1(net244),
    .X(net249));
 sky130_fd_sc_hd__mux4_4 c314 (.A0(net113),
    .A1(net207),
    .A2(net135),
    .A3(net119),
    .S0(net233),
    .S1(net920),
    .X(net250));
 sky130_fd_sc_hd__o211a_1 c315 (.A1(clknet_1_1__leaf_net130),
    .A2(net931),
    .B1(net246),
    .C1(net838),
    .X(net251));
 sky130_fd_sc_hd__or2_1 c316 (.A(net248),
    .B(net1044),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c317 (.A0(net233),
    .A1(net224),
    .A2(net215),
    .A3(net113),
    .S0(net831),
    .S1(net838),
    .X(net253));
 sky130_fd_sc_hd__and2b_2 c318 (.A_N(net122),
    .B(net819),
    .X(net254));
 sky130_fd_sc_hd__sdfstp_1 c319 (.CLK(clknet_4_7_0_clk),
    .D(net248),
    .SCD(net244),
    .SCE(net237),
    .SET_B(net819),
    .Q(net255));
 sky130_fd_sc_hd__nor3_1 c320 (.A(net923),
    .B(net955),
    .C(net831),
    .Y(net256));
 sky130_fd_sc_hd__nor3_1 c321 (.A(net118),
    .B(net239),
    .C(net838),
    .Y(net257));
 sky130_fd_sc_hd__nand3b_1 c322 (.A_N(net252),
    .B(net255),
    .C(net257),
    .Y(net258));
 sky130_fd_sc_hd__nor3_2 c323 (.A(net258),
    .B(net255),
    .C(net838),
    .Y(net985));
 sky130_fd_sc_hd__o211ai_1 c324 (.A1(net255),
    .A2(net258),
    .B1(net940),
    .C1(net213),
    .Y(net259));
 sky130_fd_sc_hd__sdfstp_1 c325 (.CLK(clknet_4_7_0_clk),
    .D(net1094),
    .SCD(net237),
    .SCE(net128),
    .SET_B(net819),
    .Q(net260));
 sky130_fd_sc_hd__sedfxbp_2 c326 (.CLK(clknet_4_12_0_clk),
    .D(net244),
    .DE(net254),
    .SCD(net985),
    .SCE(net237),
    .Q(net262),
    .Q_N(net261));
 sky130_fd_sc_hd__sedfxbp_2 c327 (.CLK(clknet_4_6_0_clk),
    .D(net259),
    .DE(net260),
    .SCD(net256),
    .SCE(net257),
    .Q(net264),
    .Q_N(net263));
 sky130_fd_sc_hd__and3b_2 c328 (.A_N(net260),
    .B(net262),
    .C(net119),
    .X(net265));
 sky130_fd_sc_hd__nor3b_1 c329 (.A(net206),
    .B(net263),
    .C_N(net831),
    .Y(net266));
 sky130_fd_sc_hd__nand3b_4 c330 (.A_N(net21),
    .B(net996),
    .C(net1023),
    .Y(net267));
 sky130_fd_sc_hd__o211ai_1 c331 (.A1(net1023),
    .A2(net1004),
    .B1(net221),
    .C1(net839),
    .Y(net268));
 sky130_fd_sc_hd__o221ai_4 c332 (.A1(net952),
    .A2(net267),
    .B1(net237),
    .B2(net220),
    .C1(net147),
    .Y(net269));
 sky130_fd_sc_hd__clkbuf_2 c333 (.A(net778),
    .X(net984));
 sky130_fd_sc_hd__o211a_4 c334 (.A1(net264),
    .A2(net267),
    .B1(clknet_1_0__leaf_net19),
    .C1(net778),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 c335 (.A(net775),
    .X(net271));
 sky130_fd_sc_hd__o211a_2 c336 (.A1(net914),
    .A2(net144),
    .B1(net267),
    .C1(clknet_1_1__leaf_net832),
    .X(net986));
 sky130_fd_sc_hd__inv_2 c337 (.A(net775),
    .Y(net272));
 sky130_fd_sc_hd__nand3_4 c338 (.A(net265),
    .B(net267),
    .C(net802),
    .Y(net273));
 sky130_fd_sc_hd__buf_6 c339 (.A(net786),
    .X(net274));
 sky130_fd_sc_hd__buf_6 c340 (.A(net778),
    .X(net275));
 sky130_fd_sc_hd__nand2_1 c341 (.A(net147),
    .B(net275),
    .Y(net276));
 sky130_fd_sc_hd__nor3b_2 c342 (.A(net144),
    .B(net115),
    .C_N(net839),
    .Y(net277));
 sky130_fd_sc_hd__and2_1 c343 (.A(net276),
    .B(net254),
    .X(net278));
 sky130_fd_sc_hd__o221a_2 c344 (.A1(net267),
    .A2(net278),
    .B1(clknet_1_1__leaf_net111),
    .B2(net952),
    .C1(net1000),
    .X(net279));
 sky130_fd_sc_hd__buf_4 c345 (.A(net776),
    .X(net280));
 sky130_fd_sc_hd__o221ai_4 c346 (.A1(net275),
    .A2(net274),
    .B1(net280),
    .B2(net794),
    .C1(net839),
    .Y(net281));
 sky130_fd_sc_hd__mux4_4 c347 (.A0(net1019),
    .A1(net275),
    .A2(net281),
    .A3(clknet_1_0__leaf_net19),
    .S0(net280),
    .S1(net802),
    .X(net282));
 sky130_fd_sc_hd__sdfbbp_1 c348 (.CLK(clknet_4_12_0_clk),
    .D(net221),
    .RESET_B(net280),
    .SCD(net1000),
    .SCE(net277),
    .SET_B(net1072),
    .Q(net284),
    .Q_N(net283));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net270),
    .A1(net280),
    .A2(net260),
    .A3(net1003),
    .S0(net283),
    .S1(net840),
    .X(net285));
 sky130_fd_sc_hd__mux4_4 c350 (.A0(clknet_1_1__leaf_net111),
    .A1(net280),
    .A2(net267),
    .A3(net960),
    .S0(net840),
    .S1(net841),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net281),
    .A1(net280),
    .A2(net1023),
    .A3(net234),
    .S0(net220),
    .S1(net778),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 c353 (.A(net804),
    .X(net991));
 sky130_fd_sc_hd__and3_1 c354 (.A(net274),
    .B(net141),
    .C(clknet_1_0__leaf_net168),
    .X(net961));
 sky130_fd_sc_hd__mux4_2 c355 (.A0(clknet_1_1__leaf_net22),
    .A1(net159),
    .A2(net1064),
    .A3(net281),
    .S0(net1019),
    .S1(net45),
    .X(net288));
 sky130_fd_sc_hd__dlymetal6s2s_1 c356 (.A(net808),
    .X(net1007));
 sky130_fd_sc_hd__o221a_4 c357 (.A1(net141),
    .A2(clknet_1_1__leaf_net175),
    .B1(clknet_1_0__leaf_net38),
    .B2(net1039),
    .C1(net842),
    .X(net289));
 sky130_fd_sc_hd__nand3b_4 c358 (.A_N(net213),
    .B(net838),
    .C(net842),
    .Y(net290));
 sky130_fd_sc_hd__o221ai_4 c359 (.A1(net290),
    .A2(net18),
    .B1(net984),
    .B2(net729),
    .C1(net842),
    .Y(net291));
 sky130_fd_sc_hd__sdfbbn_1 c360 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net168),
    .RESET_B(net291),
    .SCD(net997),
    .SCE(net159),
    .SET_B(net1019),
    .Q(net293),
    .Q_N(net292));
 sky130_fd_sc_hd__and3_4 c361 (.A(clknet_1_0__leaf_net19),
    .B(net960),
    .C(net842),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net293),
    .A1(net1009),
    .A2(net178),
    .A3(net996),
    .S0(net1004),
    .S1(net835),
    .X(net295));
 sky130_fd_sc_hd__or3_1 c363 (.A(net271),
    .B(net1044),
    .C(net42),
    .X(net296));
 sky130_fd_sc_hd__inv_1 c364 (.A(net760),
    .Y(net297));
 sky130_fd_sc_hd__nor3_1 c365 (.A(clknet_1_1__leaf_net19),
    .B(net292),
    .C(net290),
    .Y(net1010));
 sky130_fd_sc_hd__and3b_1 c366 (.A_N(net290),
    .B(net42),
    .C(net1039),
    .X(net298));
 sky130_fd_sc_hd__mux4_2 c367 (.A0(net273),
    .A1(net18),
    .A2(clknet_1_1__leaf_net169),
    .A3(net291),
    .S0(net774),
    .S1(net844),
    .X(net299));
 sky130_fd_sc_hd__o221ai_1 c368 (.A1(net298),
    .A2(net18),
    .B1(net291),
    .B2(net1019),
    .C1(clknet_1_0__leaf_net1010),
    .Y(net300));
 sky130_fd_sc_hd__mux4_2 c369 (.A0(net18),
    .A1(net1019),
    .A2(net290),
    .A3(net1044),
    .S0(clknet_1_1__leaf_net19),
    .S1(net845),
    .X(net301));
 sky130_fd_sc_hd__o221a_2 c370 (.A1(net1000),
    .A2(net291),
    .B1(clknet_1_0__leaf_net986),
    .B2(net774),
    .C1(net812),
    .X(net302));
 sky130_fd_sc_hd__inv_4 c371 (.A(net813),
    .Y(net989));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net296),
    .A1(net271),
    .A2(net178),
    .A3(clknet_1_1__leaf_net162),
    .S0(net989),
    .S1(net844),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net1007),
    .A1(net1063),
    .A2(net767),
    .A3(net842),
    .S0(net843),
    .S1(net846),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net180),
    .A1(net996),
    .A2(net1044),
    .A3(net191),
    .S0(net1007),
    .S1(net784),
    .X(net995));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net77),
    .A1(net192),
    .A2(net1014),
    .A3(net1019),
    .S0(net970),
    .S1(net960),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net58),
    .A1(net921),
    .A2(net180),
    .A3(net1019),
    .S0(net1097),
    .S1(net1080),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net291),
    .A1(net183),
    .A2(net1001),
    .A3(net989),
    .S1(net980),
    .X(net307));
 sky130_fd_sc_hd__nand2_2 c396 (.A(net957),
    .B(net201),
    .Y(net308));
 sky130_fd_sc_hd__and2_1 c397 (.A(net201),
    .B(net1021),
    .X(net309));
 sky130_fd_sc_hd__inv_4 c398 (.A(net743),
    .Y(net310));
 sky130_fd_sc_hd__buf_16 c399 (.A(net719),
    .X(net311));
 sky130_fd_sc_hd__nand2_2 c400 (.A(net210),
    .B(net199),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 c401 (.A(net719),
    .Y(net313));
 sky130_fd_sc_hd__inv_2 c402 (.A(net732),
    .Y(net314));
 sky130_fd_sc_hd__or2b_2 c403 (.A(net211),
    .B_N(net313),
    .X(net315));
 sky130_fd_sc_hd__inv_8 c404 (.A(net718),
    .Y(net316));
 sky130_fd_sc_hd__nor2_4 c405 (.A(net310),
    .B(net218),
    .Y(net317));
 sky130_fd_sc_hd__sedfxtp_4 c406 (.CLK(clknet_4_4_0_clk),
    .D(net316),
    .DE(net312),
    .SCD(net313),
    .SCE(net1015),
    .Q(net318));
 sky130_fd_sc_hd__sedfxtp_4 c407 (.CLK(clknet_4_4_0_clk),
    .D(net313),
    .DE(net317),
    .SCD(net315),
    .SCE(net1015),
    .Q(net319));
 sky130_fd_sc_hd__mux4_2 c408 (.A0(net313),
    .A1(net317),
    .A2(net199),
    .A3(net212),
    .S0(net312),
    .S1(net834),
    .X(net320));
 sky130_fd_sc_hd__or2b_1 c409 (.A(net312),
    .B_N(net317),
    .X(net321));
 sky130_fd_sc_hd__inv_6 c410 (.A(net718),
    .Y(net322));
 sky130_fd_sc_hd__mux4_1 c411 (.A0(net216),
    .A1(net321),
    .A2(net311),
    .A3(net314),
    .S0(net1033),
    .S1(net1015),
    .X(net323));
 sky130_fd_sc_hd__sedfxtp_4 c412 (.CLK(clknet_4_4_0_clk),
    .D(net311),
    .DE(net322),
    .SCD(net1033),
    .SCE(net1015),
    .Q(net324));
 sky130_fd_sc_hd__mux4_1 c413 (.A0(net321),
    .A1(net313),
    .A2(net316),
    .A3(net320),
    .S0(net317),
    .S1(net1033),
    .X(net325));
 sky130_fd_sc_hd__buf_6 c414 (.A(net746),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net314),
    .A1(net321),
    .A2(net310),
    .A3(net200),
    .S0(net1033),
    .S1(net1015),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net326),
    .A1(net324),
    .A2(net1015),
    .A3(net818),
    .S0(net990),
    .S1(net847),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net322),
    .A1(net311),
    .A2(net1041),
    .A3(net990),
    .S0(net847),
    .S1(clknet_1_1__leaf_net848),
    .X(net329));
 sky130_fd_sc_hd__o211ai_1 c418 (.A1(net74),
    .A2(net213),
    .B1(net322),
    .C1(net818),
    .Y(net330));
 sky130_fd_sc_hd__nor3_4 c419 (.A(net86),
    .B(net236),
    .C(net836),
    .Y(net994));
 sky130_fd_sc_hd__nor2b_1 c420 (.A(net226),
    .B_N(net829),
    .Y(net331));
 sky130_fd_sc_hd__nor3_1 c421 (.A(net314),
    .B(net331),
    .C(net829),
    .Y(net332));
 sky130_fd_sc_hd__buf_1 c422 (.A(net742),
    .X(net333));
 sky130_fd_sc_hd__and2b_1 c423 (.A_N(net314),
    .B(net829),
    .X(net334));
 sky130_fd_sc_hd__o221a_1 c424 (.A1(net915),
    .A2(net1030),
    .B1(net331),
    .B2(net1033),
    .C1(net1015),
    .X(net335));
 sky130_fd_sc_hd__nor2b_1 c425 (.A(net228),
    .B_N(net322),
    .Y(net336));
 sky130_fd_sc_hd__nand2b_2 c426 (.A_N(net229),
    .B(net236),
    .Y(net971));
 sky130_fd_sc_hd__clkbuf_1 c427 (.A(net742),
    .X(net337));
 sky130_fd_sc_hd__o221ai_4 c428 (.A1(net236),
    .A2(net326),
    .B1(net310),
    .B2(net739),
    .C1(net1066),
    .Y(net338));
 sky130_fd_sc_hd__mux4_1 c429 (.A0(net336),
    .A1(net1020),
    .A2(net228),
    .A3(net23),
    .S0(net1037),
    .S1(net1081),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net331),
    .A1(net229),
    .A2(net17),
    .A3(net1020),
    .S0(net994),
    .S1(net1030),
    .X(net340));
 sky130_fd_sc_hd__nand3b_2 c431 (.A_N(net927),
    .B(net450),
    .C(net739),
    .Y(net341));
 sky130_fd_sc_hd__nor3b_1 c432 (.A(net341),
    .B(net86),
    .C_N(clknet_1_1__leaf_net849),
    .Y(net342));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(clknet_1_0__leaf_net342),
    .A1(net898),
    .A2(net341),
    .A3(net330),
    .S0(net212),
    .S1(net927),
    .X(net343));
 sky130_fd_sc_hd__mux4_2 c434 (.A0(net337),
    .A1(clknet_1_0__leaf_net342),
    .A2(net994),
    .A3(net320),
    .S0(net133),
    .S1(net1066),
    .X(net344));
 sky130_fd_sc_hd__mux4_4 c435 (.A0(net1020),
    .A1(clknet_1_1__leaf_net342),
    .A2(net341),
    .A3(net739),
    .S0(net797),
    .S1(clknet_1_0__leaf_net850),
    .X(net345));
 sky130_fd_sc_hd__mux4_4 c436 (.A0(net934),
    .A1(clknet_1_1__leaf_net342),
    .A2(net92),
    .A3(net226),
    .S0(clknet_1_1__leaf_net849),
    .S1(net851),
    .X(net346));
 sky130_fd_sc_hd__mux4_2 c437 (.A0(net341),
    .A1(net1033),
    .A2(net797),
    .A3(net829),
    .S0(net851),
    .S1(net854),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net218),
    .A1(net341),
    .A2(net332),
    .A3(net347),
    .S0(clknet_1_0__leaf_net850),
    .S1(net852),
    .X(net348));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net212),
    .A1(net347),
    .A2(clknet_1_0__leaf_net342),
    .A3(clknet_1_1__leaf_net849),
    .S0(net852),
    .S1(net855),
    .X(net349));
 sky130_fd_sc_hd__or3b_1 c440 (.A(net913),
    .B(net1031),
    .C_N(net254),
    .X(net350));
 sky130_fd_sc_hd__o221a_2 c441 (.A1(net247),
    .A2(net207),
    .B1(net1030),
    .B2(net739),
    .C1(clknet_1_0__leaf_net850),
    .X(net351));
 sky130_fd_sc_hd__and3b_2 c442 (.A_N(net264),
    .B(net245),
    .C(net797),
    .X(net352));
 sky130_fd_sc_hd__sdfrbp_2 c443 (.CLK(clknet_4_6_0_clk),
    .D(net955),
    .RESET_B(net1084),
    .SCD(net1031),
    .SCE(net1018),
    .Q(net972),
    .Q_N(net353));
 sky130_fd_sc_hd__or3_1 c444 (.A(net931),
    .B(net207),
    .C(net334),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 c445 (.A(net784),
    .X(net355));
 sky130_fd_sc_hd__nand3b_2 c446 (.A_N(net355),
    .B(net354),
    .C(clknet_1_1__leaf_net850),
    .Y(net356));
 sky130_fd_sc_hd__o211ai_4 c447 (.A1(clknet_1_1__leaf_net351),
    .A2(net1031),
    .B1(net898),
    .C1(net972),
    .Y(net357));
 sky130_fd_sc_hd__nor3b_4 c448 (.A(clknet_1_0__leaf_net351),
    .B(net835),
    .C_N(clknet_1_1__leaf_net850),
    .Y(net358));
 sky130_fd_sc_hd__nand3_2 c449 (.A(net358),
    .B(net354),
    .C(net135),
    .Y(net359));
 sky130_fd_sc_hd__o211a_2 c450 (.A1(net359),
    .A2(net215),
    .B1(net355),
    .C1(net263),
    .X(net360));
 sky130_fd_sc_hd__o221ai_4 c451 (.A1(net1031),
    .A2(net319),
    .B1(net353),
    .B2(net728),
    .C1(net797),
    .Y(net361));
 sky130_fd_sc_hd__clkinv_8 c452 (.A(net784),
    .Y(net362));
 sky130_fd_sc_hd__sdfrbp_1 c453 (.CLK(clknet_4_6_0_clk),
    .D(net944),
    .RESET_B(net320),
    .SCD(net972),
    .SCE(net361),
    .Q(net987),
    .Q_N(net363));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net256),
    .A1(net119),
    .A2(net362),
    .A3(net987),
    .S0(net353),
    .S1(net856),
    .X(net364));
 sky130_fd_sc_hd__inv_4 c455 (.A(net776),
    .Y(net365));
 sky130_fd_sc_hd__buf_4 c456 (.A(net745),
    .X(net366));
 sky130_fd_sc_hd__o211ai_1 c457 (.A1(net326),
    .A2(net972),
    .B1(net1037),
    .C1(net728),
    .Y(net367));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(clknet_1_0__leaf_net351),
    .A1(net365),
    .A2(net935),
    .A3(net92),
    .S0(net364),
    .S1(net856),
    .X(net978));
 sky130_fd_sc_hd__mux4_4 c459 (.A0(net364),
    .A1(net1031),
    .A2(net898),
    .A3(net367),
    .S0(net353),
    .S1(clknet_1_0__leaf_net978),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net367),
    .A1(net366),
    .A2(net352),
    .A3(net899),
    .S0(clknet_1_1__leaf_net978),
    .S1(net853),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net135),
    .A1(clknet_1_0__leaf_net356),
    .A2(net361),
    .A3(net352),
    .S0(net365),
    .S1(net981),
    .X(net370));
 sky130_fd_sc_hd__nor3_1 c462 (.A(net365),
    .B(net334),
    .C(clknet_1_1__leaf_net832),
    .Y(net371));
 sky130_fd_sc_hd__nand3b_2 c463 (.A_N(net935),
    .B(clknet_1_0__leaf_net371),
    .C(net352),
    .Y(net372));
 sky130_fd_sc_hd__clkbuf_2 c464 (.A(net785),
    .X(net373));
 sky130_fd_sc_hd__and3b_2 c465 (.A_N(clknet_1_0__leaf_net371),
    .B(net839),
    .C(net854),
    .X(net374));
 sky130_fd_sc_hd__nor3_4 c466 (.A(net352),
    .B(net284),
    .C(net899),
    .Y(net375));
 sky130_fd_sc_hd__clkbuf_2 c467 (.A(net785),
    .X(net376));
 sky130_fd_sc_hd__o211ai_2 c468 (.A1(net149),
    .A2(net1043),
    .B1(net921),
    .C1(net920),
    .Y(net377));
 sky130_fd_sc_hd__and3_1 c469 (.A(net377),
    .B(net352),
    .C(net812),
    .X(net378));
 sky130_fd_sc_hd__or3b_1 c470 (.A(net376),
    .B(net8),
    .C_N(net260),
    .X(net379));
 sky130_fd_sc_hd__inv_1 c471 (.A(net808),
    .Y(net380));
 sky130_fd_sc_hd__clkbuf_2 c472 (.A(net800),
    .X(net381));
 sky130_fd_sc_hd__sdfbbn_1 c473 (.CLK_N(clknet_4_9_0_clk),
    .D(net373),
    .RESET_B(net381),
    .SCD(net1022),
    .SCE(net366),
    .SET_B(net365),
    .Q(net383),
    .Q_N(net382));
 sky130_fd_sc_hd__o211a_4 c474 (.A1(clknet_1_1__leaf_net371),
    .A2(net350),
    .B1(net377),
    .C1(net2),
    .X(net384));
 sky130_fd_sc_hd__inv_2 c475 (.A(net759),
    .Y(net385));
 sky130_fd_sc_hd__and3_1 c476 (.A(net385),
    .B(net261),
    .C(net818),
    .X(net386));
 sky130_fd_sc_hd__o221ai_4 c477 (.A1(net379),
    .A2(net385),
    .B1(net207),
    .B2(net8),
    .C1(net818),
    .Y(net387));
 sky130_fd_sc_hd__o221a_1 c478 (.A1(net272),
    .A2(net387),
    .B1(net381),
    .B2(net385),
    .C1(net841),
    .X(net388));
 sky130_fd_sc_hd__nor3_4 c479 (.A(net381),
    .B(net246),
    .C(net1038),
    .Y(net968));
 sky130_fd_sc_hd__sdfbbp_1 c480 (.CLK(clknet_4_9_0_clk),
    .D(net388),
    .RESET_B(net385),
    .SCD(net898),
    .SCE(net366),
    .SET_B(net1038),
    .Q(net1011),
    .Q_N(net389));
 sky130_fd_sc_hd__o221a_1 c481 (.A1(net378),
    .A2(net366),
    .B1(net365),
    .B2(net388),
    .C1(net283),
    .X(net390));
 sky130_fd_sc_hd__mux4_2 c482 (.A0(clknet_1_0__leaf_net372),
    .A1(net373),
    .A2(net388),
    .A3(net386),
    .S0(net246),
    .S1(net777),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net380),
    .A1(net373),
    .A2(net968),
    .A3(net385),
    .S0(net387),
    .S1(net840),
    .X(net392));
 sky130_fd_sc_hd__o221a_2 c484 (.A1(net171),
    .A2(net42),
    .B1(clknet_1_0__leaf_net169),
    .B2(net375),
    .C1(clknet_1_0__leaf_net34),
    .X(net393));
 sky130_fd_sc_hd__o211a_1 c485 (.A1(net334),
    .A2(net968),
    .B1(net261),
    .C1(net389),
    .X(net975));
 sky130_fd_sc_hd__o221a_4 c486 (.A1(net975),
    .A2(net1024),
    .B1(net1044),
    .B2(clknet_1_1__leaf_net303),
    .C1(net777),
    .X(net394));
 sky130_fd_sc_hd__sdfbbn_1 c487 (.CLK_N(clknet_4_9_0_clk),
    .D(net989),
    .RESET_B(clknet_1_0__leaf_net961),
    .SCD(net1024),
    .SCE(net1041),
    .SET_B(net812),
    .Q(net396),
    .Q_N(net395));
 sky130_fd_sc_hd__o221ai_4 c488 (.A1(net2),
    .A2(clknet_1_0__leaf_net304),
    .B1(net375),
    .B2(net395),
    .C1(clknet_1_1__leaf_net303),
    .Y(net397));
 sky130_fd_sc_hd__sdfrtn_1 c489 (.CLK_N(clknet_4_11_0_clk),
    .D(net375),
    .RESET_B(net1068),
    .SCD(clknet_1_0__leaf_net34),
    .SCE(net843),
    .Q(net979));
 sky130_fd_sc_hd__mux4_4 c490 (.A0(net396),
    .A1(net988),
    .A2(net979),
    .A3(net170),
    .S0(net375),
    .S1(clknet_1_1__leaf_net34),
    .X(net398));
 sky130_fd_sc_hd__o221a_1 c491 (.A1(net322),
    .A2(net968),
    .B1(net979),
    .B2(net899),
    .C1(clknet_1_0__leaf_net34),
    .X(net399));
 sky130_fd_sc_hd__o221a_4 c492 (.A1(net159),
    .A2(net273),
    .B1(clknet_1_1__leaf_net169),
    .B2(net170),
    .C1(net823),
    .X(net400));
 sky130_fd_sc_hd__sdfbbn_1 c493 (.CLK_N(clknet_4_9_0_clk),
    .D(net375),
    .RESET_B(clknet_1_1__leaf_net372),
    .SCD(net395),
    .SCE(net985),
    .SET_B(net823),
    .Q(net976),
    .Q_N(net401));
 sky130_fd_sc_hd__sdfbbp_1 c494 (.CLK(clknet_4_11_0_clk),
    .D(net991),
    .RESET_B(net401),
    .SCD(net392),
    .SCE(net964),
    .SET_B(net1076),
    .Q(net403),
    .Q_N(net402));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net262),
    .A1(net281),
    .A2(net941),
    .A3(net899),
    .S0(net401),
    .S1(net809),
    .X(net404));
 sky130_fd_sc_hd__mux4_4 c496 (.A0(net404),
    .A1(net1062),
    .A2(net976),
    .A3(net402),
    .S0(clknet_1_0__leaf_net162),
    .S1(net988),
    .X(net405));
 sky130_fd_sc_hd__mux4_4 c497 (.A0(net403),
    .A1(net1041),
    .A2(clknet_1_1__leaf_net1008),
    .A3(net41),
    .S0(net401),
    .S1(net977),
    .X(net406));
 sky130_fd_sc_hd__mux4_4 c498 (.A0(net392),
    .A1(net213),
    .A2(net403),
    .A3(net171),
    .S0(clknet_1_0__leaf_net304),
    .S1(net985),
    .X(net407));
 sky130_fd_sc_hd__mux4_2 c499 (.A0(net366),
    .A1(net991),
    .A2(net403),
    .A3(clknet_1_0__leaf_net961),
    .S0(net159),
    .S1(clknet_1_0__leaf_net34),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net402),
    .A1(net1043),
    .A2(net71),
    .A3(net979),
    .S0(net815),
    .S1(net859),
    .X(net409));
 sky130_fd_sc_hd__sdfbbn_1 c501 (.CLK_N(clknet_4_11_0_clk),
    .D(net71),
    .RESET_B(net2),
    .SCD(net1087),
    .SCE(net159),
    .SET_B(net1088),
    .Q(net411),
    .Q_N(net410));
 sky130_fd_sc_hd__mux4_2 c502 (.A0(clknet_1_1__leaf_net304),
    .A1(net410),
    .A2(net366),
    .A3(clknet_1_1__leaf_net303),
    .S0(net784),
    .S1(net859),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net411),
    .A1(net409),
    .A2(net401),
    .A3(net809),
    .S0(net859),
    .S1(net860),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net413),
    .A1(net411),
    .A2(net979),
    .A3(net941),
    .S0(net859),
    .S1(net860),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net899),
    .A1(net409),
    .A2(net404),
    .A3(net976),
    .S0(net375),
    .S1(net410),
    .X(net415));
 sky130_fd_sc_hd__buf_4 c528 (.A(net733),
    .X(net416));
 sky130_fd_sc_hd__and2_4 c529 (.A(net329),
    .B(net990),
    .X(net417));
 sky130_fd_sc_hd__nor2_2 c530 (.A(net416),
    .B(clknet_1_0__leaf_net848),
    .Y(net418));
 sky130_fd_sc_hd__inv_1 c531 (.A(net733),
    .Y(net419));
 sky130_fd_sc_hd__inv_4 c532 (.A(net776),
    .Y(net420));
 sky130_fd_sc_hd__and2_1 c533 (.A(net943),
    .B(net420),
    .X(net421));
 sky130_fd_sc_hd__nand2b_4 c534 (.A_N(net420),
    .B(net416),
    .Y(net422));
 sky130_fd_sc_hd__nor3_2 c535 (.A(net419),
    .B(net1033),
    .C(net422),
    .Y(net423));
 sky130_fd_sc_hd__o211ai_4 c536 (.A1(net421),
    .A2(net422),
    .B1(net423),
    .C1(net1043),
    .Y(net424));
 sky130_fd_sc_hd__or2_2 c537 (.A(net420),
    .B(clknet_1_0__leaf_net418),
    .X(net425));
 sky130_fd_sc_hd__and2_1 c538 (.A(net423),
    .B(net421),
    .X(net426));
 sky130_fd_sc_hd__or2_2 c539 (.A(net1043),
    .B(clknet_1_0__leaf_net418),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 c540 (.A(net732),
    .X(net428));
 sky130_fd_sc_hd__and2_0 c541 (.A(net92),
    .B(clknet_1_0__leaf_net418),
    .X(net429));
 sky130_fd_sc_hd__and2_0 c542 (.A(net428),
    .B(clknet_1_0__leaf_net425),
    .X(net430));
 sky130_fd_sc_hd__buf_1 c543 (.A(net792),
    .X(net431));
 sky130_fd_sc_hd__nor3_2 c544 (.A(net431),
    .B(net199),
    .C(clknet_1_1__leaf_net418),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 c545 (.A(net807),
    .Y(net433));
 sky130_fd_sc_hd__clkbuf_2 c546 (.A(net1089),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(net434),
    .A1(net422),
    .A2(net419),
    .A3(net421),
    .S0(net424),
    .S1(clknet_1_0__leaf_net429),
    .X(net435));
 sky130_fd_sc_hd__sdfbbn_1 c548 (.CLK_N(clknet_4_1_0_clk),
    .D(clknet_1_1__leaf_net425),
    .RESET_B(net426),
    .SCD(net308),
    .SCE(clknet_1_0__leaf_net429),
    .SET_B(net861),
    .Q(net437),
    .Q_N(net436));
 sky130_fd_sc_hd__nand3_1 c549 (.A(clknet_1_1__leaf_net432),
    .B(net437),
    .C(net861),
    .Y(net438));
 sky130_fd_sc_hd__or2_1 c550 (.A(net318),
    .B(net847),
    .X(net439));
 sky130_fd_sc_hd__and2_1 c551 (.A(net436),
    .B(net818),
    .X(net440));
 sky130_fd_sc_hd__inv_4 c552 (.A(net773),
    .Y(net441));
 sky130_fd_sc_hd__clkbuf_1 c553 (.A(net773),
    .X(net442));
 sky130_fd_sc_hd__nor2_1 c554 (.A(net439),
    .B(net1081),
    .Y(net443));
 sky130_fd_sc_hd__o221a_4 c555 (.A1(net441),
    .A2(net310),
    .B1(net1037),
    .B2(clknet_1_0__leaf_net427),
    .C1(net436),
    .X(net444));
 sky130_fd_sc_hd__o211a_4 c556 (.A1(net440),
    .A2(clknet_1_1__leaf_net427),
    .B1(net570),
    .C1(net836),
    .X(net445));
 sky130_fd_sc_hd__nor2_2 c557 (.A(net152),
    .B(net440),
    .Y(net446));
 sky130_fd_sc_hd__sdfbbp_1 c558 (.CLK(clknet_4_1_0_clk),
    .D(net443),
    .RESET_B(net338),
    .SCD(clknet_1_0__leaf_net445),
    .SCE(net923),
    .SET_B(clknet_1_0__leaf_net849),
    .Q(net448),
    .Q_N(net447));
 sky130_fd_sc_hd__or2b_1 c559 (.A(net338),
    .B_N(net852),
    .X(net449));
 sky130_fd_sc_hd__inv_12 c695_12 (.A(clknet_1_0__leaf_net967),
    .Y(net1057));
 sky130_fd_sc_hd__and3b_1 c561 (.A_N(net1033),
    .B(net1030),
    .C(net837),
    .X(net451));
 sky130_fd_sc_hd__nand2b_1 c562 (.A_N(net437),
    .B(net442),
    .Y(net452));
 sky130_fd_sc_hd__inv_6 c563 (.A(net801),
    .Y(net453));
 sky130_fd_sc_hd__buf_6 c564 (.A(net807),
    .X(net454));
 sky130_fd_sc_hd__and3_1 c565 (.A(net452),
    .B(net449),
    .C(net433),
    .X(net455));
 sky130_fd_sc_hd__o211a_1 c566 (.A1(net448),
    .A2(net455),
    .B1(net433),
    .C1(net861),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 c567 (.A(net801),
    .X(net457));
 sky130_fd_sc_hd__or3_4 c568 (.A(net433),
    .B(net453),
    .C(net1028),
    .X(net458));
 sky130_fd_sc_hd__sdfbbn_2 c569 (.CLK_N(clknet_4_1_0_clk),
    .D(net316),
    .RESET_B(net447),
    .SCD(net458),
    .SCE(clknet_1_1__leaf_net445),
    .SET_B(net1027),
    .Q(net460),
    .Q_N(net459));
 sky130_fd_sc_hd__o211ai_1 c570 (.A1(net1027),
    .A2(net455),
    .B1(net459),
    .C1(net752),
    .Y(net461));
 sky130_fd_sc_hd__sdfbbn_1 c571 (.CLK_N(clknet_4_1_0_clk),
    .D(net455),
    .RESET_B(net454),
    .SCD(clknet_1_1__leaf_net427),
    .SCE(net1028),
    .SET_B(net752),
    .Q(net463),
    .Q_N(net462));
 sky130_fd_sc_hd__nand3_4 c572 (.A(net460),
    .B(clknet_1_1__leaf_net429),
    .C(net1030),
    .Y(net464));
 sky130_fd_sc_hd__o221ai_4 c573 (.A1(net940),
    .A2(net460),
    .B1(clknet_1_1__leaf_net429),
    .B2(clknet_1_1__leaf_net417),
    .C1(net362),
    .Y(net465));
 sky130_fd_sc_hd__o221a_2 c574 (.A1(net362),
    .A2(clknet_1_1__leaf_net429),
    .B1(net1020),
    .B2(net1037),
    .C1(net1030),
    .X(net466));
 sky130_fd_sc_hd__inv_1 c575 (.A(net1090),
    .Y(net467));
 sky130_fd_sc_hd__clkbuf_2 c576 (.A(net786),
    .X(net468));
 sky130_fd_sc_hd__o221a_1 c577 (.A1(net460),
    .A2(net468),
    .B1(net711),
    .B2(net799),
    .C1(net857),
    .X(net469));
 sky130_fd_sc_hd__o221a_1 c578 (.A1(net308),
    .A2(net318),
    .B1(net446),
    .B2(net857),
    .C1(net862),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 c579 (.A(net800),
    .X(net471));
 sky130_fd_sc_hd__mux4_2 c580 (.A0(net469),
    .A1(net1040),
    .A2(clknet_1_1__leaf_net445),
    .A3(clknet_1_1__leaf_net417),
    .S0(net1020),
    .S1(net1030),
    .X(net472));
 sky130_fd_sc_hd__inv_2 c581 (.A(net776),
    .Y(net473));
 sky130_fd_sc_hd__mux4_2 c582 (.A0(net473),
    .A1(clknet_1_0__leaf_net417),
    .A2(net469),
    .A3(net921),
    .S0(net940),
    .S1(net862),
    .X(net474));
 sky130_fd_sc_hd__mux4_4 c583 (.A0(net470),
    .A1(net1037),
    .A2(clknet_1_0__leaf_net429),
    .A3(net728),
    .S0(net863),
    .S1(net865),
    .X(net475));
 sky130_fd_sc_hd__o221ai_4 c584 (.A1(net950),
    .A2(net318),
    .B1(net446),
    .B2(net857),
    .C1(net865),
    .Y(net476));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net469),
    .A1(net1030),
    .A2(net476),
    .A3(net857),
    .S0(net862),
    .S1(net865),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net1037),
    .A1(net927),
    .A2(net463),
    .A3(net800),
    .S0(net864),
    .S1(net865),
    .X(net478));
 sky130_fd_sc_hd__sdfbbp_1 c587 (.CLK(clknet_4_3_0_clk),
    .D(net467),
    .RESET_B(net362),
    .SCD(net476),
    .SCE(net857),
    .SET_B(net1074),
    .Q(net480),
    .Q_N(net479));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net478),
    .A1(net480),
    .A2(net125),
    .A3(net254),
    .S0(net459),
    .S1(net1028),
    .X(net481));
 sky130_fd_sc_hd__mux4_4 c589 (.A0(net468),
    .A1(net478),
    .A2(net1037),
    .A3(net481),
    .S0(net981),
    .S1(net865),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(clknet_1_1__leaf_net429),
    .A1(net481),
    .A2(net468),
    .A3(net476),
    .S0(net799),
    .S1(net867),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net446),
    .A1(net480),
    .A2(net972),
    .A3(net468),
    .S0(net1028),
    .S1(net862),
    .X(net484));
 sky130_fd_sc_hd__mux4_4 c592 (.A0(net247),
    .A1(net478),
    .A2(net479),
    .A3(clknet_1_1__leaf_net429),
    .S0(net800),
    .S1(net866),
    .X(net485));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net471),
    .A1(net463),
    .A2(clknet_1_1__leaf_net485),
    .A3(clknet_1_1__leaf_net417),
    .S0(net468),
    .S1(net712),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_2 c594 (.A(net814),
    .X(net487));
 sky130_fd_sc_hd__o211a_1 c595 (.A1(net422),
    .A2(net1038),
    .B1(net1029),
    .C1(net841),
    .X(net488));
 sky130_fd_sc_hd__o221a_1 c596 (.A1(net386),
    .A2(net260),
    .B1(net1022),
    .B2(net207),
    .C1(net484),
    .X(net489));
 sky130_fd_sc_hd__mux4_4 c597 (.A0(net264),
    .A1(net1020),
    .A2(net353),
    .A3(net1045),
    .S0(clknet_1_0__leaf_net464),
    .S1(net1037),
    .X(net490));
 sky130_fd_sc_hd__o221a_2 c598 (.A1(net1045),
    .A2(net376),
    .B1(net476),
    .B2(net1038),
    .C1(clknet_1_0__leaf_net832),
    .X(net491));
 sky130_fd_sc_hd__o221ai_1 c599 (.A1(net207),
    .A2(net8),
    .B1(net1033),
    .B2(net840),
    .C1(clknet_1_0__leaf_net869),
    .Y(net492));
 sky130_fd_sc_hd__mux4_4 c600 (.A0(net422),
    .A1(net283),
    .A2(clknet_1_0__leaf_net372),
    .A3(net712),
    .S0(clknet_1_1__leaf_net992),
    .S1(clknet_1_0__leaf_net868),
    .X(net493));
 sky130_fd_sc_hd__sdfbbn_1 c601 (.CLK_N(clknet_4_9_0_clk),
    .D(net484),
    .RESET_B(net1029),
    .SCD(net476),
    .SCE(net1038),
    .SET_B(net1022),
    .Q(net495),
    .Q_N(net494));
 sky130_fd_sc_hd__o221a_4 c602 (.A1(net492),
    .A2(net142),
    .B1(net1029),
    .B2(net990),
    .C1(clknet_1_0__leaf_net868),
    .X(net496));
 sky130_fd_sc_hd__sdfbbn_1 c603 (.CLK_N(clknet_4_9_0_clk),
    .D(net1022),
    .RESET_B(net1020),
    .SCD(net422),
    .SCE(net1040),
    .SET_B(clknet_1_1__leaf_net869),
    .Q(net498),
    .Q_N(net497));
 sky130_fd_sc_hd__o221a_2 c604 (.A1(net476),
    .A2(net277),
    .B1(net281),
    .B2(clknet_1_0__leaf_net496),
    .C1(clknet_1_0__leaf_net969),
    .X(net499));
 sky130_fd_sc_hd__o221ai_4 c605 (.A1(net487),
    .A2(net8),
    .B1(net981),
    .B2(net866),
    .C1(clknet_1_0__leaf_net969),
    .Y(net500));
 sky130_fd_sc_hd__o221a_1 c606 (.A1(net487),
    .A2(net498),
    .B1(net494),
    .B2(net1020),
    .C1(net1012),
    .X(net501));
 sky130_fd_sc_hd__o221a_1 c607 (.A1(net246),
    .A2(net500),
    .B1(net386),
    .B2(net320),
    .C1(clknet_1_0__leaf_net832),
    .X(net502));
 sky130_fd_sc_hd__or3b_1 c608 (.A(net497),
    .B(clknet_1_1__leaf_net967),
    .C_N(net1013),
    .X(net503));
 sky130_fd_sc_hd__o221ai_1 c609 (.A1(net385),
    .A2(net387),
    .B1(net487),
    .B2(clknet_1_1__leaf_net503),
    .C1(clknet_1_0__leaf_net869),
    .Y(net504));
 sky130_fd_sc_hd__mux4_4 c610 (.A0(net488),
    .A1(clknet_1_0__leaf_net503),
    .A2(net497),
    .A3(clknet_1_0__leaf_net504),
    .S0(net1029),
    .S1(net811),
    .X(net505));
 sky130_fd_sc_hd__mux4_2 c611 (.A0(net495),
    .A1(clknet_1_0__leaf_net503),
    .A2(net284),
    .A3(clknet_1_1__leaf_net504),
    .S0(net1040),
    .S1(net92),
    .X(net506));
 sky130_fd_sc_hd__mux4_4 c612 (.A0(net387),
    .A1(net495),
    .A2(clknet_1_0__leaf_net504),
    .A3(clknet_1_0__leaf_net503),
    .S0(net811),
    .S1(net870),
    .X(net507));
 sky130_fd_sc_hd__buf_2 c613 (.A(net814),
    .X(net508));
 sky130_fd_sc_hd__mux4_2 c614 (.A0(clknet_1_1__leaf_net496),
    .A1(clknet_1_1__leaf_net503),
    .A2(net142),
    .A3(net353),
    .S0(net494),
    .S1(net870),
    .X(net509));
 sky130_fd_sc_hd__mux4_2 c615 (.A0(net509),
    .A1(net495),
    .A2(net488),
    .A3(clknet_1_0__leaf_net503),
    .S0(net508),
    .S1(net963),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net262),
    .A1(clknet_1_0__leaf_net34),
    .A2(net971),
    .A3(net846),
    .S0(net981),
    .S1(net873),
    .X(net511));
 sky130_fd_sc_hd__mux4_4 c617 (.A0(clknet_1_0__leaf_net169),
    .A1(net972),
    .A2(net320),
    .A3(net858),
    .S0(net1032),
    .S1(clknet_1_1__leaf_net868),
    .X(net512));
 sky130_fd_sc_hd__mux4_2 c618 (.A0(net281),
    .A1(net1038),
    .A2(net1040),
    .A3(net1045),
    .S0(net844),
    .S1(net867),
    .X(net513));
 sky130_fd_sc_hd__mux4_4 c619 (.A0(net498),
    .A1(net1011),
    .A2(clknet_1_0__leaf_net162),
    .A3(clknet_1_1__leaf_net464),
    .S0(net835),
    .S1(net1032),
    .X(net514));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net945),
    .A1(net951),
    .A2(net939),
    .A3(net937),
    .S0(net3),
    .S1(net1044),
    .X(net0));
 sky130_fd_sc_hd__mux4_2 c620 (.A0(clknet_1_0__leaf_net303),
    .A1(net513),
    .A2(net498),
    .A3(net1029),
    .S0(net1032),
    .S1(net875),
    .X(net515));
 sky130_fd_sc_hd__mux4_4 c621 (.A0(clknet_1_0__leaf_net162),
    .A1(net923),
    .A2(net1061),
    .A3(net1024),
    .S0(net840),
    .S1(net981),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(clknet_1_0__leaf_net34),
    .A1(clknet_1_0__leaf_net303),
    .A2(net780),
    .A3(net960),
    .S0(net843),
    .S1(net1032),
    .X(net517));
 sky130_fd_sc_hd__mux4_2 c623 (.A0(net320),
    .A1(net513),
    .A2(clknet_1_0__leaf_net464),
    .A3(net963),
    .S0(clknet_1_1__leaf_net992),
    .S1(clknet_1_1__leaf_net868),
    .X(net518));
 sky130_fd_sc_hd__mux4_4 c624 (.A0(net1043),
    .A1(clknet_1_1__leaf_net372),
    .A2(net1011),
    .A3(net1038),
    .S0(net422),
    .S1(net870),
    .X(net519));
 sky130_fd_sc_hd__mux4_4 c625 (.A0(net1038),
    .A1(clknet_1_1__leaf_net516),
    .A2(net968),
    .A3(net389),
    .S0(net840),
    .S1(net858),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net513),
    .A1(net389),
    .A2(net796),
    .A3(net825),
    .S0(net858),
    .S1(net874),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net927),
    .A1(net487),
    .A2(net1024),
    .A3(net1040),
    .S0(net972),
    .S1(net977),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net522),
    .A1(net42),
    .A2(clknet_1_0__leaf_net961),
    .A3(net1029),
    .S0(net844),
    .S1(net990),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net521),
    .A1(net1024),
    .A2(net513),
    .A3(clknet_1_0__leaf_net162),
    .S0(net816),
    .S1(net1032),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c63 (.A0(net946),
    .A1(net938),
    .A2(net948),
    .A3(net942),
    .S0(net3),
    .S1(net939),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(clknet_1_0__leaf_net34),
    .A1(net521),
    .A2(clknet_1_0__leaf_net169),
    .A3(net825),
    .S0(net1032),
    .S1(net973),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net422),
    .A1(net293),
    .A2(net513),
    .A3(net968),
    .S0(net780),
    .S1(net858),
    .X(net965));
 sky130_fd_sc_hd__mux4_2 c632 (.A0(net965),
    .A1(clknet_1_1__leaf_net464),
    .A2(net513),
    .A3(net508),
    .S0(net803),
    .S1(net815),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net1029),
    .A1(net521),
    .A2(net422),
    .A3(net513),
    .S0(net845),
    .S1(net867),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net1024),
    .A1(net42),
    .A2(net835),
    .A3(net1032),
    .S0(net867),
    .S1(net876),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net528),
    .A1(net1029),
    .A2(clknet_1_0__leaf_net169),
    .A3(net422),
    .S0(clknet_1_1__leaf_net969),
    .S1(net876),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net1060),
    .A1(net528),
    .A2(net41),
    .A3(net816),
    .S0(net990),
    .S1(net877),
    .X(net530));
 sky130_fd_sc_hd__mux4_4 c637 (.A0(net530),
    .A1(net284),
    .A2(net920),
    .A3(net971),
    .S0(net840),
    .S1(net877),
    .X(net531));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net952),
    .A1(net950),
    .A2(net956),
    .A3(net3),
    .S0(net0),
    .S1(net939),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net928),
    .A1(net914),
    .A2(net919),
    .A3(net912),
    .S0(net900),
    .S1(net913),
    .X(net3));
 sky130_fd_sc_hd__nand2_1 c66 (.A(net931),
    .B(net1045),
    .Y(net4));
 sky130_fd_sc_hd__or2b_4 c660 (.A(net81),
    .B_N(net434),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_1 c661 (.A(net806),
    .X(net533));
 sky130_fd_sc_hd__inv_2 c662 (.A(net646),
    .Y(net534));
 sky130_fd_sc_hd__buf_16 c663 (.A(net645),
    .X(net535));
 sky130_fd_sc_hd__nand3_1 c664 (.A(clknet_1_0__leaf_net432),
    .B(net215),
    .C(net81),
    .Y(net536));
 sky130_fd_sc_hd__inv_4 c665 (.A(net817),
    .Y(net537));
 sky130_fd_sc_hd__sdfrtp_2 c666 (.CLK(clknet_4_0_0_clk),
    .D(net424),
    .RESET_B(net532),
    .SCD(net78),
    .SCE(net1026),
    .Q(net538));
 sky130_fd_sc_hd__inv_6 c667 (.A(net817),
    .Y(net539));
 sky130_fd_sc_hd__inv_1 c668 (.A(net761),
    .Y(net540));
 sky130_fd_sc_hd__nand2b_1 c669 (.A_N(net86),
    .B(clknet_1_0__leaf_net848),
    .Y(net541));
 sky130_fd_sc_hd__nor3b_4 c67 (.A(net951),
    .B(net1044),
    .C_N(net0),
    .Y(net5));
 sky130_fd_sc_hd__or2_1 c670 (.A(net540),
    .B(net204),
    .X(net542));
 sky130_fd_sc_hd__or2_2 c671 (.A(net416),
    .B(net542),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c672 (.A0(clknet_1_0__leaf_net536),
    .A1(clknet_1_0__leaf_net541),
    .A2(net317),
    .A3(net534),
    .S0(net539),
    .S1(net1016),
    .X(net544));
 sky130_fd_sc_hd__buf_6 c673 (.A(net792),
    .X(net545));
 sky130_fd_sc_hd__nand2b_1 c674 (.A_N(clknet_1_1__leaf_net541),
    .B(net545),
    .Y(net546));
 sky130_fd_sc_hd__nand2_1 c675 (.A(net317),
    .B(net204),
    .Y(net547));
 sky130_fd_sc_hd__mux4_2 c676 (.A0(net533),
    .A1(net543),
    .A2(net539),
    .A3(net540),
    .S0(net545),
    .S1(net879),
    .X(net548));
 sky130_fd_sc_hd__inv_2 c677 (.A(net1077),
    .Y(net549));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net208),
    .A1(net542),
    .A2(net549),
    .A3(net548),
    .S0(net1069),
    .S1(net1067),
    .X(net550));
 sky130_fd_sc_hd__or3_4 c679 (.A(net545),
    .B(net543),
    .C(net772),
    .X(net551));
 sky130_fd_sc_hd__and2_1 c68 (.A(net927),
    .B(net917),
    .X(net6));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(net549),
    .A1(net551),
    .A2(net317),
    .A3(net548),
    .S0(net532),
    .S1(net543),
    .X(net552));
 sky130_fd_sc_hd__sdfbbp_1 c681 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_1__leaf_net438),
    .RESET_B(net548),
    .SCD(net551),
    .SCE(net324),
    .SET_B(net1078),
    .Q(net554),
    .Q_N(net553));
 sky130_fd_sc_hd__nand3b_1 c682 (.A_N(net537),
    .B(net547),
    .C(net1040),
    .Y(net555));
 sky130_fd_sc_hd__sdfrtp_4 c683 (.CLK(clknet_4_0_0_clk),
    .D(net548),
    .RESET_B(net1067),
    .SCD(net1027),
    .SCE(net879),
    .Q(net556));
 sky130_fd_sc_hd__o211a_1 c684 (.A1(net554),
    .A2(net1026),
    .B1(net1045),
    .C1(net879),
    .X(net557));
 sky130_fd_sc_hd__nand3_2 c685 (.A(net557),
    .B(net537),
    .C(net556),
    .Y(net558));
 sky130_fd_sc_hd__o211a_1 c686 (.A1(net558),
    .A2(net547),
    .B1(net548),
    .C1(net1027),
    .X(net559));
 sky130_fd_sc_hd__sdfbbn_1 c687 (.CLK_N(clknet_4_0_0_clk),
    .D(net543),
    .RESET_B(net558),
    .SCD(net78),
    .SCE(net555),
    .SET_B(net553),
    .Q(net561),
    .Q_N(net560));
 sky130_fd_sc_hd__sdfrtp_4 c688 (.CLK(clknet_4_0_0_clk),
    .D(net555),
    .RESET_B(net1069),
    .SCD(net557),
    .SCE(net1027),
    .Q(net562));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net547),
    .A1(net555),
    .A2(net556),
    .A3(net543),
    .S0(net561),
    .S1(net1026),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 c69 (.A(net661),
    .X(net7));
 sky130_fd_sc_hd__sdfbbn_2 c690 (.CLK_N(clknet_4_0_0_clk),
    .D(net200),
    .RESET_B(net558),
    .SCD(net1045),
    .SCE(net557),
    .SET_B(net556),
    .Q(net565),
    .Q_N(net564));
 sky130_fd_sc_hd__mux4_4 c691 (.A0(net85),
    .A1(net558),
    .A2(net545),
    .A3(net557),
    .S0(net458),
    .S1(net880),
    .X(net566));
 sky130_fd_sc_hd__o221a_1 c692 (.A1(net454),
    .A2(net554),
    .B1(net564),
    .B2(net458),
    .C1(net1027),
    .X(net567));
 sky130_fd_sc_hd__o221ai_1 c693 (.A1(net567),
    .A2(net448),
    .B1(net562),
    .B2(net537),
    .C1(net1027),
    .Y(net568));
 sky130_fd_sc_hd__mux4_4 c694 (.A0(net561),
    .A1(net538),
    .A2(net1043),
    .A3(net556),
    .S0(net85),
    .S1(net1027),
    .X(net569));
 sky130_fd_sc_hd__clkinv_2 c352_13 (.A(net804),
    .Y(net1058));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net569),
    .A1(net923),
    .A2(net553),
    .A3(net564),
    .S0(net454),
    .S1(net560),
    .X(net571));
 sky130_fd_sc_hd__and3b_1 c697 (.A_N(net538),
    .B(net556),
    .C(net458),
    .X(net572));
 sky130_fd_sc_hd__o221a_2 c698 (.A1(net1057),
    .A2(net548),
    .B1(net572),
    .B2(net560),
    .C1(net1026),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net566),
    .A1(net458),
    .A2(net556),
    .A3(net1026),
    .S0(net564),
    .S1(net883),
    .X(net574));
 sky130_fd_sc_hd__inv_6 c70 (.A(net661),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net572),
    .A1(net557),
    .A2(net556),
    .A3(net454),
    .S0(net1027),
    .S1(net795),
    .X(net575));
 sky130_fd_sc_hd__sdfbbp_1 c701 (.CLK(clknet_4_0_0_clk),
    .D(net1091),
    .RESET_B(net1069),
    .SCD(net532),
    .SCE(net572),
    .SET_B(net1027),
    .Q(net577),
    .Q_N(net576));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net575),
    .A1(net577),
    .A2(net558),
    .A3(net538),
    .S0(net572),
    .S1(net761),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net78),
    .A1(net562),
    .A2(net572),
    .A3(net577),
    .S0(net564),
    .S1(net883),
    .X(net579));
 sky130_fd_sc_hd__sdfbbn_2 c704 (.CLK_N(clknet_4_2_0_clk),
    .D(clknet_1_0__leaf_net485),
    .RESET_B(net1092),
    .SCD(net577),
    .SCE(net562),
    .SET_B(net882),
    .Q(net581),
    .Q_N(net580));
 sky130_fd_sc_hd__o221a_4 c705 (.A1(net318),
    .A2(net125),
    .B1(net565),
    .B2(clknet_1_1__leaf_net485),
    .C1(net1026),
    .X(net582));
 sky130_fd_sc_hd__mux4_4 c706 (.A0(clknet_1_1__leaf_net485),
    .A1(net1026),
    .A2(net581),
    .A3(net458),
    .S0(net994),
    .S1(net864),
    .X(net583));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_4_2_0_clk),
    .D(net577),
    .RESET_B(clknet_1_0__leaf_net546),
    .SCD(net458),
    .SCE(net580),
    .SET_B(net880),
    .Q(net585),
    .Q_N(net584));
 sky130_fd_sc_hd__o211a_1 c708 (.A1(net1026),
    .A2(net125),
    .B1(net921),
    .C1(net864),
    .X(net586));
 sky130_fd_sc_hd__o221ai_1 c709 (.A1(net565),
    .A2(net920),
    .B1(net580),
    .B2(net1037),
    .C1(net883),
    .Y(net587));
 sky130_fd_sc_hd__or2b_2 c71 (.A(net7),
    .B_N(net900),
    .X(net9));
 sky130_fd_sc_hd__o221ai_4 c710 (.A1(net585),
    .A2(net921),
    .B1(net1043),
    .B2(net1037),
    .C1(net817),
    .Y(net588));
 sky130_fd_sc_hd__o221a_1 c711 (.A1(net215),
    .A2(net1026),
    .B1(net576),
    .B2(net866),
    .C1(net882),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(clknet_1_0__leaf_net546),
    .A1(net589),
    .A2(net577),
    .A3(net584),
    .S0(net1028),
    .S1(net728),
    .X(net590));
 sky130_fd_sc_hd__o211ai_1 c713 (.A1(net585),
    .A2(net125),
    .B1(net589),
    .C1(net883),
    .Y(net591));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net589),
    .A1(net579),
    .A2(net1040),
    .A3(net580),
    .S0(net532),
    .S1(net882),
    .X(net592));
 sky130_fd_sc_hd__o221ai_1 c715 (.A1(net576),
    .A2(net761),
    .B1(net817),
    .B2(net866),
    .C1(net1095),
    .Y(net593));
 sky130_fd_sc_hd__sdfbbp_1 c716 (.CLK(clknet_4_2_0_clk),
    .D(net593),
    .RESET_B(clknet_1_0__leaf_net485),
    .SCD(net535),
    .SCE(net580),
    .SET_B(net863),
    .Q(net595),
    .Q_N(net594));
 sky130_fd_sc_hd__o221a_1 c717 (.A1(net458),
    .A2(net584),
    .B1(net565),
    .B2(net588),
    .C1(net576),
    .X(net596));
 sky130_fd_sc_hd__sdfbbn_1 c718 (.CLK_N(clknet_4_3_0_clk),
    .D(net532),
    .RESET_B(net595),
    .SCD(net565),
    .SCE(net863),
    .SET_B(net881),
    .Q(net598),
    .Q_N(net597));
 sky130_fd_sc_hd__mux4_2 c719 (.A0(net586),
    .A1(net125),
    .A2(net576),
    .A3(net458),
    .S0(net588),
    .S1(net885),
    .X(net599));
 sky130_fd_sc_hd__o211a_1 c72 (.A1(net8),
    .A2(net1022),
    .B1(net952),
    .C1(net1),
    .X(net10));
 sky130_fd_sc_hd__mux4_4 c720 (.A0(net596),
    .A1(net599),
    .A2(net458),
    .A3(net795),
    .S0(net882),
    .S1(net885),
    .X(net600));
 sky130_fd_sc_hd__o221ai_4 c721 (.A1(net586),
    .A2(net594),
    .B1(net867),
    .B2(net883),
    .C1(net886),
    .Y(net601));
 sky130_fd_sc_hd__o221a_1 c722 (.A1(net581),
    .A2(clknet_1_0__leaf_net485),
    .B1(net601),
    .B2(net125),
    .C1(net758),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net599),
    .A1(net581),
    .A2(net1043),
    .A3(net758),
    .S0(net885),
    .S1(net1093),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net601),
    .A1(net599),
    .A2(net589),
    .A3(net597),
    .S0(net923),
    .S1(net795),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net587),
    .A1(net596),
    .A2(net565),
    .A3(net758),
    .S0(net795),
    .S1(net886),
    .X(net605));
 sky130_fd_sc_hd__mux4_4 c726 (.A0(net581),
    .A1(net1017),
    .A2(net923),
    .A3(net866),
    .S0(net871),
    .S1(net873),
    .X(net606));
 sky130_fd_sc_hd__o221ai_1 c727 (.A1(net142),
    .A2(net588),
    .B1(net562),
    .B2(net551),
    .C1(net886),
    .Y(net607));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net254),
    .A1(net376),
    .A2(net551),
    .A3(net8),
    .S0(net791),
    .S1(net884),
    .X(net608));
 sky130_fd_sc_hd__mux4_4 c729 (.A0(net1017),
    .A1(net551),
    .A2(net580),
    .A3(net8),
    .S0(net866),
    .S1(net871),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_4 c73 (.A(net669),
    .X(net11));
 sky130_fd_sc_hd__mux4_4 c730 (.A0(net551),
    .A1(net598),
    .A2(net562),
    .A3(net799),
    .S0(clknet_1_0__leaf_net832),
    .S1(clknet_1_1__leaf_net992),
    .X(net610));
 sky130_fd_sc_hd__mux4_4 c731 (.A0(net599),
    .A1(net284),
    .A2(net562),
    .A3(net921),
    .S0(clknet_1_0__leaf_net868),
    .S1(clknet_1_0__leaf_net888),
    .X(net611));
 sky130_fd_sc_hd__mux4_2 c732 (.A0(net382),
    .A1(net1043),
    .A2(net283),
    .A3(net791),
    .S0(net798),
    .S1(clknet_1_0__leaf_net887),
    .X(net612));
 sky130_fd_sc_hd__mux4_2 c733 (.A0(clknet_1_1__leaf_net374),
    .A1(net595),
    .A2(net8),
    .A3(net1017),
    .S0(net1029),
    .S1(net866),
    .X(net613));
 sky130_fd_sc_hd__mux4_2 c734 (.A0(clknet_1_0__leaf_net612),
    .A1(clknet_1_0__leaf_net374),
    .A2(net283),
    .A3(net921),
    .S0(net885),
    .S1(clknet_1_0__leaf_net888),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net601),
    .A1(clknet_1_0__leaf_net546),
    .A2(net581),
    .A3(net1045),
    .S0(clknet_1_0__leaf_net992),
    .S1(net881),
    .X(net615));
 sky130_fd_sc_hd__o221a_2 c736 (.A1(net581),
    .A2(net383),
    .B1(clknet_1_1__leaf_net612),
    .B2(net798),
    .C1(net811),
    .X(net616));
 sky130_fd_sc_hd__mux4_4 c737 (.A0(clknet_1_1__leaf_net616),
    .A1(net376),
    .A2(net254),
    .A3(clknet_1_0__leaf_net770),
    .S0(net821),
    .S1(net881),
    .X(net617));
 sky130_fd_sc_hd__o221ai_2 c738 (.A1(net8),
    .A2(net921),
    .B1(net562),
    .B2(net551),
    .C1(net811),
    .Y(net618));
 sky130_fd_sc_hd__mux4_2 c739 (.A0(net387),
    .A1(clknet_1_0__leaf_net464),
    .A2(clknet_1_1__leaf_net617),
    .A3(net142),
    .S0(net803),
    .S1(net884),
    .X(net619));
 sky130_fd_sc_hd__buf_16 c74 (.A(clknet_1_0__leaf_net769),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net383),
    .A1(net125),
    .A2(net1017),
    .A3(clknet_1_0__leaf_net616),
    .S0(net1038),
    .S1(clknet_1_0__leaf_net868),
    .X(net620));
 sky130_fd_sc_hd__mux4_4 c741 (.A0(clknet_1_1__leaf_net617),
    .A1(net824),
    .A2(net963),
    .A3(clknet_1_0__leaf_net832),
    .S0(clknet_1_0__leaf_net868),
    .S1(net890),
    .X(net621));
 sky130_fd_sc_hd__o221ai_4 c742 (.A1(net562),
    .A2(net601),
    .B1(clknet_1_0__leaf_net374),
    .B2(clknet_1_1__leaf_net888),
    .C1(net891),
    .Y(net622));
 sky130_fd_sc_hd__o221ai_4 c743 (.A1(clknet_1_0__leaf_net617),
    .A2(net1017),
    .B1(net822),
    .B2(net880),
    .C1(net890),
    .Y(net623));
 sky130_fd_sc_hd__o221a_2 c744 (.A1(clknet_1_0__leaf_net617),
    .A2(net1017),
    .B1(clknet_1_1__leaf_net616),
    .B2(net822),
    .C1(net881),
    .X(net624));
 sky130_fd_sc_hd__mux4_4 c745 (.A0(net142),
    .A1(clknet_1_0__leaf_net612),
    .A2(clknet_1_0__leaf_net617),
    .A3(clknet_1_0__leaf_net546),
    .S0(net821),
    .S1(clknet_1_0__leaf_net889),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(clknet_1_0__leaf_net616),
    .A1(net920),
    .A2(clknet_1_1__leaf_net464),
    .A3(clknet_1_1__leaf_net770),
    .S0(net796),
    .S1(net890),
    .X(net626));
 sky130_fd_sc_hd__mux4_4 c747 (.A0(clknet_1_1__leaf_net617),
    .A1(net508),
    .A2(net387),
    .A3(net785),
    .S0(net880),
    .S1(net892),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net72),
    .A1(net1045),
    .A2(net866),
    .A3(net873),
    .S0(net875),
    .S1(net894),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net284),
    .A1(net923),
    .A2(clknet_1_0__leaf_net992),
    .A3(net874),
    .S0(clknet_1_1__leaf_net889),
    .S1(net891),
    .X(net629));
 sky130_fd_sc_hd__inv_8 c75 (.A(net788),
    .Y(net13));
 sky130_fd_sc_hd__mux4_4 c750 (.A0(clknet_1_1__leaf_net546),
    .A1(net867),
    .A2(net871),
    .A3(net872),
    .S0(net891),
    .S1(net893),
    .X(net630));
 sky130_fd_sc_hd__mux4_4 c751 (.A0(net1045),
    .A1(net799),
    .A2(net874),
    .A3(net878),
    .S0(net892),
    .S1(net895),
    .X(net631));
 sky130_fd_sc_hd__mux4_2 c752 (.A0(net588),
    .A1(clknet_1_0__leaf_net992),
    .A2(net878),
    .A3(clknet_1_1__leaf_net889),
    .S0(net891),
    .S1(net895),
    .X(net632));
 sky130_fd_sc_hd__mux4_2 c753 (.A0(net628),
    .A1(net632),
    .A2(net588),
    .A3(net867),
    .S0(net874),
    .S1(net893),
    .X(net633));
 sky130_fd_sc_hd__mux4_4 c754 (.A0(net631),
    .A1(net923),
    .A2(net781),
    .A3(clknet_1_1__leaf_net992),
    .S0(net875),
    .S1(net894),
    .X(net634));
 sky130_fd_sc_hd__mux4_2 c755 (.A0(net588),
    .A1(clknet_1_0__leaf_net516),
    .A2(net508),
    .A3(net796),
    .S0(clknet_1_1__leaf_net868),
    .S1(net894),
    .X(net635));
 sky130_fd_sc_hd__mux4_4 c756 (.A0(net72),
    .A1(net283),
    .A2(net796),
    .A3(net866),
    .S0(net878),
    .S1(net896),
    .X(net636));
 sky130_fd_sc_hd__mux4_4 c757 (.A0(clknet_1_1__leaf_net464),
    .A1(net906),
    .A2(clknet_1_1__leaf_net546),
    .A3(net781),
    .S0(clknet_1_1__leaf_net887),
    .S1(net896),
    .X(net637));
 sky130_fd_sc_hd__mux4_2 c758 (.A0(net629),
    .A1(net866),
    .A2(clknet_1_1__leaf_net868),
    .A3(net894),
    .S0(net896),
    .S1(net897),
    .X(net638));
 sky130_fd_sc_hd__mux4_2 c759 (.A0(net508),
    .A1(clknet_1_1__leaf_net464),
    .A2(clknet_1_0__leaf_net887),
    .A3(clknet_1_0__leaf_net889),
    .S0(net895),
    .S1(net896),
    .X(net639));
 sky130_fd_sc_hd__o211a_2 c76 (.A1(net6),
    .A2(net4),
    .B1(net11),
    .C1(net13),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net636),
    .A1(clknet_1_1__leaf_net546),
    .A2(net872),
    .A3(clknet_1_1__leaf_net887),
    .S0(net896),
    .S1(net897),
    .X(net640));
 sky130_fd_sc_hd__mux4_2 c761 (.A0(net598),
    .A1(net824),
    .A2(net871),
    .A3(clknet_1_1__leaf_net889),
    .S0(net896),
    .S1(net897),
    .X(net641));
 sky130_fd_sc_hd__mux4_4 c762 (.A0(net634),
    .A1(net284),
    .A2(clknet_1_1__leaf_net546),
    .A3(net867),
    .S0(net893),
    .S1(net896),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net641),
    .A1(net508),
    .A2(net803),
    .A3(net875),
    .S0(net884),
    .S1(net896),
    .X(net643));
 sky130_fd_sc_hd__mux4_2 c764 (.A0(net638),
    .A1(net643),
    .A2(net508),
    .A3(net803),
    .S0(net875),
    .S1(net895));
 sky130_fd_sc_hd__mux4_1 c77 (.A0(net6),
    .A1(net924),
    .A2(net926),
    .A3(clknet_1_0__leaf_net12),
    .S0(net1022),
    .S1(net3),
    .X(net15));
 sky130_fd_sc_hd__o211a_2 c78 (.A1(clknet_1_0__leaf_net12),
    .A2(net14),
    .B1(net949),
    .C1(net926),
    .X(net16));
 sky130_fd_sc_hd__inv_4 c85_8 (.A(net771),
    .Y(net1053));
 sky130_fd_sc_hd__clkinv_8 c80 (.A(net669),
    .Y(net18));
 sky130_fd_sc_hd__and3b_1 c81 (.A_N(net9),
    .B(net1051),
    .C(net740),
    .X(net19));
 sky130_fd_sc_hd__or2b_1 c82 (.A(net920),
    .B_N(net740),
    .X(net20));
 sky130_fd_sc_hd__clkinv_4 c83 (.A(net790),
    .Y(net21));
 sky130_fd_sc_hd__or3_4 c84 (.A(net1050),
    .B(net912),
    .C(clknet_1_0__leaf_net12),
    .X(net22));
 sky130_fd_sc_hd__clkinv_4 c560_11 (.A(clknet_1_1__leaf_net967),
    .Y(net1056));
 sky130_fd_sc_hd__o211ai_4 c86 (.A1(net21),
    .A2(net1054),
    .B1(net20),
    .C1(net11),
    .Y(net24));
 sky130_fd_sc_hd__o211ai_4 c87 (.A1(clknet_1_0__leaf_net24),
    .A2(net1053),
    .B1(clknet_1_0__leaf_net22),
    .C1(net21),
    .Y(net25));
 sky130_fd_sc_hd__nand2_2 c88 (.A(net4),
    .B(net14),
    .Y(net982));
 sky130_fd_sc_hd__inv_6 c89 (.A(net760),
    .Y(net26));
 sky130_fd_sc_hd__nor2_1 c90 (.A(net13),
    .B(net947),
    .Y(net27));
 sky130_fd_sc_hd__buf_2 c91 (.A(net760),
    .X(net28));
 sky130_fd_sc_hd__nor2_4 c92 (.A(net1049),
    .B(net27),
    .Y(net29));
 sky130_fd_sc_hd__or3_2 c93 (.A(net7),
    .B(net13),
    .C(clknet_1_0__leaf_net29),
    .X(net30));
 sky130_fd_sc_hd__nand2b_1 c94 (.A_N(net27),
    .B(net953),
    .Y(net31));
 sky130_fd_sc_hd__or2_1 c95 (.A(net946),
    .B(net927),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 c96 (.A(net805),
    .X(net33));
 sky130_fd_sc_hd__nor2_2 c97 (.A(clknet_1_1__leaf_net29),
    .B(net26),
    .Y(net34));
 sky130_fd_sc_hd__nand2b_1 c98 (.A_N(net32),
    .B(net33),
    .Y(net35));
 sky130_fd_sc_hd__or2b_2 c99 (.A(net33),
    .B_N(net928),
    .X(net36));
 sky130_fd_sc_hd__mux4_1 merge765 (.A0(net332),
    .A1(net200),
    .A2(net308),
    .A3(net330),
    .S0(net336),
    .S1(net1030),
    .X(net644));
 sky130_fd_sc_hd__sdfsbp_1 merge766 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net430),
    .SCD(clknet_1_0__leaf_net438),
    .SCE(net204),
    .SET_B(net532),
    .Q(net646),
    .Q_N(net645));
 sky130_fd_sc_hd__o221ai_1 merge767 (.A1(net930),
    .A2(net80),
    .B1(net102),
    .B2(net95),
    .C1(net1035),
    .Y(net647));
 sky130_fd_sc_hd__o211ai_1 merge768 (.A1(net103),
    .A2(net122),
    .B1(net124),
    .C1(net121),
    .Y(net648));
 sky130_fd_sc_hd__o211a_1 merge769 (.A1(net76),
    .A2(net1040),
    .B1(net909),
    .C1(net80),
    .X(net649));
 sky130_fd_sc_hd__o211a_1 merge770 (.A1(net200),
    .A2(net81),
    .B1(net205),
    .C1(net203),
    .X(net650));
 sky130_fd_sc_hd__o211ai_1 merge771 (.A1(net0),
    .A2(net1004),
    .B1(net234),
    .C1(net267),
    .Y(net651));
 sky130_fd_sc_hd__o211ai_1 merge772 (.A1(net223),
    .A2(net224),
    .B1(net205),
    .C1(net233),
    .Y(net652));
 sky130_fd_sc_hd__o221a_1 merge773 (.A1(net1030),
    .A2(clknet_1_1__leaf_net445),
    .B1(clknet_1_0__leaf_net417),
    .B2(net362),
    .C1(net861),
    .X(net653));
 sky130_fd_sc_hd__inv_4 merge774 (.A(net777),
    .Y(net654));
 sky130_fd_sc_hd__o221ai_2 merge775 (.A1(net239),
    .A2(net234),
    .B1(net128),
    .B2(net237),
    .C1(clknet_1_0__leaf_net130),
    .Y(net655));
 sky130_fd_sc_hd__mux4_2 merge776 (.A0(net1033),
    .A1(net476),
    .A2(net246),
    .A3(clknet_1_1__leaf_net504),
    .S0(net494),
    .S1(clknet_1_1__leaf_net503),
    .X(net656));
 sky130_fd_sc_hd__o211a_1 merge777 (.A1(net928),
    .A2(net1014),
    .B1(net26),
    .C1(clknet_1_1__leaf_net25),
    .X(net657));
 sky130_fd_sc_hd__o211ai_1 merge778 (.A1(net347),
    .A2(clknet_1_1__leaf_net427),
    .B1(clknet_1_0__leaf_net849),
    .C1(net851),
    .Y(net658));
 sky130_fd_sc_hd__o211ai_2 merge779 (.A1(net91),
    .A2(net315),
    .B1(clknet_1_0__leaf_net417),
    .C1(net316),
    .Y(net659));
 sky130_fd_sc_hd__o211ai_1 merge780 (.A1(net90),
    .A2(net898),
    .B1(net308),
    .C1(net1015),
    .Y(net660));
 sky130_fd_sc_hd__inv_2 merge781 (.A(net793),
    .Y(net661));
 sky130_fd_sc_hd__mux4_2 merge782 (.A0(net18),
    .A1(net1004),
    .A2(net55),
    .A3(net912),
    .S0(clknet_1_1__leaf_net160),
    .S1(net779),
    .X(net662));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(clknet_1_1__leaf_net356),
    .A1(net363),
    .A2(net277),
    .A3(net350),
    .S0(net281),
    .S1(net835),
    .X(net663));
 sky130_fd_sc_hd__o211a_1 merge784 (.A1(net1047),
    .A2(net1000),
    .B1(clknet_1_0__leaf_net167),
    .C1(net729),
    .X(net664));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net354),
    .A1(net1018),
    .A2(clknet_1_1__leaf_net351),
    .A3(net357),
    .S0(net333),
    .S1(net839),
    .X(net665));
 sky130_fd_sc_hd__mux4_1 merge786 (.A0(net278),
    .A1(clknet_1_1__leaf_net34),
    .A2(net45),
    .A3(net178),
    .S0(net1059),
    .S1(net1019),
    .X(net666));
 sky130_fd_sc_hd__o211a_2 merge787 (.A1(clknet_1_1__leaf_net111),
    .A2(net146),
    .B1(net1003),
    .C1(net820),
    .X(net667));
 sky130_fd_sc_hd__o221ai_2 merge788 (.A1(clknet_1_0__leaf_net16),
    .A2(net0),
    .B1(net224),
    .B2(net21),
    .C1(net1000),
    .Y(net668));
 sky130_fd_sc_hd__clkinv_4 merge789 (.A(net810),
    .Y(net669));
 sky130_fd_sc_hd__mux4_4 merge790 (.A0(net568),
    .A1(net562),
    .A2(net454),
    .A3(net442),
    .S0(clknet_1_0__leaf_net445),
    .S1(net1020),
    .X(net670));
 sky130_fd_sc_hd__o211ai_4 merge791 (.A1(net315),
    .A2(clknet_1_0__leaf_net427),
    .B1(net76),
    .C1(net1016),
    .Y(net671));
 sky130_fd_sc_hd__mux4_2 merge792 (.A0(clknet_1_1__leaf_net372),
    .A1(net1022),
    .A2(net988),
    .A3(clknet_1_0__leaf_net175),
    .S0(net150),
    .S1(net1075),
    .X(net672));
 sky130_fd_sc_hd__o211ai_4 merge793 (.A1(net434),
    .A2(net1016),
    .B1(clknet_1_0__leaf_net438),
    .C1(net424),
    .Y(net673));
 sky130_fd_sc_hd__mux4_4 merge794 (.A0(net297),
    .A1(net273),
    .A2(clknet_1_1__leaf_net34),
    .A3(net127),
    .S0(net1000),
    .S1(net1065),
    .X(net674));
 sky130_fd_sc_hd__mux4_4 merge795 (.A0(net948),
    .A1(net1003),
    .A2(clknet_1_0__leaf_net1008),
    .A3(net294),
    .S0(net290),
    .S1(clknet_1_0__leaf_net961),
    .X(net675));
 sky130_fd_sc_hd__o211a_1 merge796 (.A1(net213),
    .A2(net209),
    .B1(net238),
    .C1(net234),
    .X(net676));
 sky130_fd_sc_hd__o211a_1 merge797 (.A1(net315),
    .A2(net1015),
    .B1(net320),
    .C1(net1082),
    .X(net677));
 sky130_fd_sc_hd__o211ai_1 merge798 (.A1(net206),
    .A2(net203),
    .B1(net80),
    .C1(net958),
    .Y(net678));
 sky130_fd_sc_hd__o211ai_1 merge799 (.A1(net237),
    .A2(net73),
    .B1(net200),
    .C1(net812),
    .Y(net679));
 sky130_fd_sc_hd__o221ai_1 merge800 (.A1(net539),
    .A2(clknet_1_1__leaf_net536),
    .B1(net534),
    .B2(net548),
    .C1(net547),
    .Y(net680));
 sky130_fd_sc_hd__mux4_2 merge801 (.A0(net13),
    .A1(clknet_1_1__leaf_net16),
    .A2(net8),
    .A3(net95),
    .S0(net103),
    .S1(net102),
    .X(net681));
 sky130_fd_sc_hd__mux4_2 merge802 (.A0(net245),
    .A1(clknet_1_0__leaf_net464),
    .A2(clknet_1_1__leaf_net429),
    .A3(net361),
    .S0(net1041),
    .S1(net990),
    .X(net682));
 sky130_fd_sc_hd__mux4_1 merge803 (.A0(net119),
    .A1(net361),
    .A2(net353),
    .A3(net88),
    .S0(net124),
    .S1(net114),
    .X(net683));
 sky130_fd_sc_hd__mux4_2 merge804 (.A0(clknet_1_1__leaf_net110),
    .A1(net106),
    .A2(net96),
    .A3(net273),
    .S0(net213),
    .S1(net818),
    .X(net684));
 sky130_fd_sc_hd__o211ai_4 merge805 (.A1(clknet_1_1__leaf_net38),
    .A2(net982),
    .B1(net65),
    .C1(net826),
    .Y(net685));
 sky130_fd_sc_hd__mux4_1 merge806 (.A0(clknet_1_1__leaf_net30),
    .A1(net26),
    .A2(net11),
    .A3(net182),
    .S0(net180),
    .S1(net1005),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 merge807 (.A0(net1),
    .A1(net11),
    .A2(net1022),
    .A3(net937),
    .S0(net126),
    .S1(net121),
    .X(net687));
 sky130_fd_sc_hd__mux4_4 merge808 (.A0(net898),
    .A1(net320),
    .A2(net277),
    .A3(net462),
    .S0(clknet_1_1__leaf_net417),
    .S1(net468),
    .X(net688));
 sky130_fd_sc_hd__mux4_4 merge809 (.A0(net230),
    .A1(net234),
    .A2(net78),
    .A3(net114),
    .S0(net265),
    .S1(net237),
    .X(net689));
 sky130_fd_sc_hd__o221ai_4 merge810 (.A1(net129),
    .A2(net147),
    .B1(net5),
    .B2(net9),
    .C1(net952),
    .Y(net690));
 sky130_fd_sc_hd__mux4_1 merge811 (.A0(net81),
    .A1(net87),
    .A2(net201),
    .A3(net203),
    .S0(net202),
    .S1(net763),
    .X(net691));
 sky130_fd_sc_hd__o221a_1 merge812 (.A1(net121),
    .A2(net900),
    .B1(net952),
    .B2(net123),
    .C1(net128),
    .X(net692));
 sky130_fd_sc_hd__mux4_2 merge813 (.A0(net96),
    .A1(net142),
    .A2(clknet_1_1__leaf_net16),
    .A3(net4),
    .S0(clknet_1_0__leaf_net19),
    .S1(net5),
    .X(net693));
 sky130_fd_sc_hd__mux4_1 merge814 (.A0(net324),
    .A1(net311),
    .A2(net1015),
    .A3(net907),
    .S0(net200),
    .S1(net204),
    .X(net694));
 sky130_fd_sc_hd__mux4_1 merge815 (.A0(net11),
    .A1(clknet_1_0__leaf_net16),
    .A2(clknet_1_0__leaf_net22),
    .A3(net151),
    .S0(clknet_1_0__leaf_net140),
    .S1(net136),
    .X(net695));
 sky130_fd_sc_hd__mux4_1 merge816 (.A0(net203),
    .A1(net199),
    .A2(net200),
    .A3(net945),
    .S0(net233),
    .S1(net914),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 merge817 (.A0(net82),
    .A1(net317),
    .A2(net1016),
    .A3(net237),
    .S0(net220),
    .S1(net1022),
    .X(net697));
 sky130_fd_sc_hd__mux4_1 merge818 (.A0(clknet_1_1__leaf_net418),
    .A1(net1056),
    .A2(net200),
    .A3(net455),
    .S0(net453),
    .S1(net454),
    .X(net698));
 sky130_fd_sc_hd__mux4_1 merge819 (.A0(net1014),
    .A1(net1001),
    .A2(net5),
    .A3(net6),
    .S0(net900),
    .S1(net813),
    .X(net699));
 sky130_fd_sc_hd__mux4_1 merge820 (.A0(net423),
    .A1(net424),
    .A2(clknet_1_0__leaf_net429),
    .A3(net542),
    .S0(net1026),
    .S1(net532),
    .X(net700));
 sky130_fd_sc_hd__mux4_1 merge821 (.A0(net919),
    .A1(net80),
    .A2(net143),
    .A3(net11),
    .S0(net1014),
    .S1(net1025),
    .X(net701));
 sky130_fd_sc_hd__mux4_1 merge822 (.A0(net199),
    .A1(net1016),
    .A2(net146),
    .A3(net148),
    .S0(net1000),
    .S1(net833),
    .X(net702));
 sky130_fd_sc_hd__o221a_1 merge823 (.A1(net87),
    .A2(net205),
    .B1(net203),
    .B2(net1021),
    .C1(net912),
    .X(net703));
 sky130_fd_sc_hd__mux4_1 merge824 (.A0(clknet_1_0__leaf_net427),
    .A1(net426),
    .A2(clknet_1_1__leaf_net432),
    .A3(net451),
    .S0(net444),
    .S1(net449),
    .X(net704));
 sky130_fd_sc_hd__mux4_2 merge825 (.A0(net426),
    .A1(clknet_1_0__leaf_net432),
    .A2(net428),
    .A3(net86),
    .S0(net324),
    .S1(clknet_1_1__leaf_net430),
    .X(net705));
 sky130_fd_sc_hd__mux4_2 merge826 (.A0(net900),
    .A1(net1042),
    .A2(net1014),
    .A3(clknet_1_1__leaf_net140),
    .S0(net1039),
    .S1(clknet_1_0__leaf_net25),
    .X(net706));
 sky130_fd_sc_hd__mux4_4 merge827 (.A0(net80),
    .A1(net136),
    .A2(net902),
    .A3(net5),
    .S0(clknet_1_1__leaf_net16),
    .S1(net740),
    .X(net707));
 sky130_fd_sc_hd__and2b_1 merge828 (.A_N(net456),
    .B(net461),
    .X(net708));
 sky130_fd_sc_hd__nand2b_1 merge829 (.A_N(net649),
    .B(net691),
    .Y(net709));
 sky130_fd_sc_hd__or2_1 merge830 (.A(net117),
    .B(net104),
    .X(net710));
 sky130_fd_sc_hd__dfrbp_1 merge831 (.CLK(clknet_4_3_0_clk),
    .D(net483),
    .RESET_B(net465),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__and2_4 merge832 (.A(net300),
    .B(net301),
    .X(net713));
 sky130_fd_sc_hd__and2b_2 merge833 (.A_N(net489),
    .B(net491),
    .X(net714));
 sky130_fd_sc_hd__nand2_4 merge834 (.A(net269),
    .B(net286),
    .Y(net715));
 sky130_fd_sc_hd__and2_2 merge835 (.A(net390),
    .B(net391),
    .X(net716));
 sky130_fd_sc_hd__or2_4 merge836 (.A(net630),
    .B(net633),
    .X(net717));
 sky130_fd_sc_hd__dfrbp_2 merge837 (.CLK(clknet_4_4_0_clk),
    .D(net660),
    .RESET_B(net677),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__nand2b_2 merge838 (.A_N(net590),
    .B(net602),
    .Y(net720));
 sky130_fd_sc_hd__dfrtn_1 merge839 (.CLK_N(clknet_4_13_0_clk),
    .D(net154),
    .RESET_B(net667),
    .Q(net721));
 sky130_fd_sc_hd__nand2b_2 merge840 (.A_N(net186),
    .B(net189),
    .Y(net722));
 sky130_fd_sc_hd__and2_2 merge841 (.A(net559),
    .B(net573),
    .X(net723));
 sky130_fd_sc_hd__nor2_4 merge842 (.A(net515),
    .B(net519),
    .Y(net724));
 sky130_fd_sc_hd__dfrtp_1 merge843 (.CLK(clknet_4_13_0_clk),
    .RESET_B(net44),
    .Q(net46));
 sky130_fd_sc_hd__or2b_1 merge844 (.A(net225),
    .B_N(net240),
    .X(net726));
 sky130_fd_sc_hd__nor2b_1 merge845 (.A(net552),
    .B_N(net550),
    .Y(net727));
 sky130_fd_sc_hd__dfrtp_4 merge846 (.CLK(clknet_4_6_0_clk),
    .D(net360),
    .RESET_B(net370),
    .Q(net728));
 sky130_fd_sc_hd__dfrtp_4 merge847 (.CLK(clknet_4_13_0_clk),
    .D(net158),
    .RESET_B(net165),
    .Q(net729));
 sky130_fd_sc_hd__or2_1 merge848 (.A(net606),
    .B(net607),
    .X(net730));
 sky130_fd_sc_hd__nand2b_1 merge849 (.A_N(net393),
    .B(net394),
    .Y(net731));
 sky130_fd_sc_hd__dfsbp_1 merge850 (.CLK(clknet_4_1_0_clk),
    .D(net659),
    .SET_B(net671),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__dfsbp_1 merge851 (.CLK(clknet_4_5_0_clk),
    .D(net650),
    .SET_B(net676),
    .Q(net735),
    .Q_N(net734));
 sky130_fd_sc_hd__nand2_1 merge852 (.A(net138),
    .B(net648),
    .Y(net736));
 sky130_fd_sc_hd__nor2_1 merge853 (.A(net251),
    .B(net249),
    .Y(net737));
 sky130_fd_sc_hd__nor2_4 merge854 (.A(net57),
    .B(net66),
    .Y(net738));
 sky130_fd_sc_hd__dfstp_2 merge855 (.CLK(clknet_4_4_0_clk),
    .D(net335),
    .SET_B(net339),
    .Q(net739));
 sky130_fd_sc_hd__dfstp_1 merge856 (.CLK(clknet_4_13_0_clk),
    .D(net10),
    .SET_B(net15),
    .Q(net740));
 sky130_fd_sc_hd__dfstp_1 merge857 (.CLK(clknet_4_14_0_clk),
    .SET_B(net306),
    .Q(net307));
 sky130_fd_sc_hd__nor2b_1 merge858 (.A(net198),
    .B_N(net407),
    .Y(net741));
 sky130_fd_sc_hd__dlrbn_2 merge859 (.D(net702),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net644),
    .Q(net743),
    .Q_N(net742));
 sky130_fd_sc_hd__and2b_2 merge860 (.A_N(net197),
    .B(net194),
    .X(net744));
 sky130_fd_sc_hd__dlrbn_2 merge861 (.D(net694),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net683),
    .Q(net746),
    .Q_N(net745));
 sky130_fd_sc_hd__and2b_1 merge862 (.A_N(net287),
    .B(net713),
    .X(net747));
 sky130_fd_sc_hd__dlrbp_2 merge863 (.D(net678),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net696),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__or2_1 merge864 (.A(net618),
    .B(net642),
    .X(net750));
 sky130_fd_sc_hd__dlrbp_2 merge865 (.D(net708),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net703),
    .Q(net752),
    .Q_N(net751));
 sky130_fd_sc_hd__nor2b_1 merge866 (.A(net574),
    .B_N(net578),
    .Y(net753));
 sky130_fd_sc_hd__and2b_1 merge867 (.A_N(net525),
    .B(net640),
    .X(net754));
 sky130_fd_sc_hd__and2b_4 merge868 (.A_N(net400),
    .B(net415),
    .X(net755));
 sky130_fd_sc_hd__or2b_4 merge869 (.A(net608),
    .B_N(net639),
    .X(net756));
 sky130_fd_sc_hd__and2b_1 merge870 (.A_N(net501),
    .B(net527),
    .X(net757));
 sky130_fd_sc_hd__dlrtn_1 merge871 (.D(net604),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net720),
    .Q(net758));
 sky130_fd_sc_hd__dlrtn_2 merge872 (.D(net647),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net684),
    .Q(net759));
 sky130_fd_sc_hd__dlrtn_2 merge873 (.D(net657),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net675),
    .Q(net760));
 sky130_fd_sc_hd__dlrtp_2 merge874 (.D(net680),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net723),
    .Q(net761));
 sky130_fd_sc_hd__or2_1 merge875 (.A(net619),
    .B(net506),
    .X(net762));
 sky130_fd_sc_hd__dlrtp_2 merge876 (.D(net692),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net84),
    .Q(net763));
 sky130_fd_sc_hd__nand2b_1 merge877 (.A_N(net399),
    .B(net523),
    .Y(net764));
 sky130_fd_sc_hd__dlrtp_4 merge878 (.D(net710),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net709),
    .Q(net765));
 sky130_fd_sc_hd__nor2_4 merge879 (.A(net520),
    .B(net625),
    .Y(net766));
 sky130_fd_sc_hd__edfxbp_1 merge880 (.CLK(clknet_4_14_0_clk),
    .D(net193),
    .DE(net302),
    .Q(net999),
    .Q_N(net767));
 sky130_fd_sc_hd__edfxtp_1 merge881 (.CLK(clknet_4_7_0_clk),
    .D(net652),
    .DE(net655),
    .Q(net768));
 sky130_fd_sc_hd__sdlclkp_1 merge882 (.CLK(clknet_4_13_0_clk),
    .GATE(net166),
    .SCE(net687),
    .GCLK(net769));
 sky130_fd_sc_hd__sdlclkp_2 merge883 (.CLK(clknet_4_8_0_clk),
    .GATE(net611),
    .SCE(net624),
    .GCLK(net770));
 sky130_fd_sc_hd__sdlclkp_4 merge884 (.CLK(clknet_4_13_0_clk),
    .GATE(net681),
    .SCE(net695),
    .GCLK(net771));
 sky130_fd_sc_hd__dfrbp_1 merge885 (.CLK(clknet_4_1_0_clk),
    .D(net658),
    .RESET_B(net727),
    .Q(net773),
    .Q_N(net772));
 sky130_fd_sc_hd__dfrbp_1 merge886 (.CLK(clknet_4_14_0_clk),
    .D(net755),
    .RESET_B(net289),
    .Q(net964),
    .Q_N(net774));
 sky130_fd_sc_hd__dfrtn_1 merge887 (.CLK_N(clknet_4_6_0_clk),
    .D(net651),
    .RESET_B(net679),
    .Q(net775));
 sky130_fd_sc_hd__dfrtp_4 merge888 (.CLK(clknet_4_6_0_clk),
    .D(net697),
    .RESET_B(net682),
    .Q(net776));
 sky130_fd_sc_hd__dfrtp_4 merge889 (.CLK(clknet_4_9_0_clk),
    .D(net716),
    .RESET_B(net701),
    .Q(net777));
 sky130_fd_sc_hd__dfrtp_2 merge890 (.CLK(clknet_4_12_0_clk),
    .D(net715),
    .RESET_B(net668),
    .Q(net778));
 sky130_fd_sc_hd__dfsbp_1 merge891 (.CLK(clknet_4_15_0_clk),
    .D(net177),
    .SET_B(net744),
    .Q(net779),
    .Q_N(net1005));
 sky130_fd_sc_hd__dfsbp_1 merge892 (.CLK(clknet_4_11_0_clk),
    .D(net511),
    .SET_B(net514),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__nand2_4 merge893 (.A(net613),
    .B(net623),
    .Y(net782));
 sky130_fd_sc_hd__nor2_1 merge894 (.A(net622),
    .B(net615),
    .Y(net783));
 sky130_fd_sc_hd__dfstp_4 merge895 (.CLK(clknet_4_12_0_clk),
    .D(net665),
    .SET_B(net741),
    .Q(net784));
 sky130_fd_sc_hd__dfstp_1 merge896 (.CLK(clknet_4_8_0_clk),
    .D(net621),
    .SET_B(net663),
    .Q(net785));
 sky130_fd_sc_hd__dfstp_2 merge897 (.CLK(clknet_4_6_0_clk),
    .D(net653),
    .SET_B(net689),
    .Q(net786));
 sky130_fd_sc_hd__dlrbn_2 merge898 (.D(net690),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net722),
    .Q(net788),
    .Q_N(net787));
 sky130_fd_sc_hd__dlrbn_2 merge899 (.D(net693),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net706),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dlrbp_1 merge900 (.D(net700),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net605),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dlrbp_1 merge901 (.D(net279),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net699),
    .Q(net794),
    .Q_N(net793));
 sky130_fd_sc_hd__dlrtn_1 merge902 (.D(net753),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net603),
    .Q(net795));
 sky130_fd_sc_hd__dlrtn_1 merge903 (.D(net717),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net766),
    .Q(net796));
 sky130_fd_sc_hd__dlrtn_2 merge904 (.D(net349),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net344),
    .Q(net797));
 sky130_fd_sc_hd__dlrtp_2 merge905 (.D(net730),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net662),
    .Q(net798));
 sky130_fd_sc_hd__dlrtp_1 merge906 (.D(net466),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net591),
    .Q(net799));
 sky130_fd_sc_hd__dlrtp_1 merge907 (.D(net477),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net688),
    .Q(net800));
 sky130_fd_sc_hd__edfxbp_1 merge908 (.CLK(clknet_4_3_0_clk),
    .D(net268),
    .DE(net698),
    .Q(net802),
    .Q_N(net801));
 sky130_fd_sc_hd__edfxtp_1 merge909 (.CLK(clknet_4_10_0_clk),
    .D(net750),
    .DE(net754),
    .Q(net803));
 sky130_fd_sc_hd__sdlclkp_1 merge910 (.CLK(clknet_4_3_0_clk),
    .GATE(net757),
    .SCE(net670),
    .GCLK(net967));
 sky130_fd_sc_hd__sdlclkp_2 merge911 (.CLK(clknet_4_14_0_clk),
    .GATE(net666),
    .SCE(net664),
    .GCLK(net804));
 sky130_fd_sc_hd__sdlclkp_4 merge912 (.CLK(clknet_4_15_0_clk),
    .GATE(net686),
    .SCE(net196),
    .GCLK(net805));
 sky130_fd_sc_hd__dfrbp_1 merge913 (.CLK(clknet_4_1_0_clk),
    .D(net704),
    .RESET_B(net705),
    .Q(net807),
    .Q_N(net806));
 sky130_fd_sc_hd__dfrbp_1 merge914 (.CLK(clknet_4_9_0_clk),
    .D(net397),
    .RESET_B(net672),
    .Q(net809),
    .Q_N(net808));
 sky130_fd_sc_hd__dfrtn_1 merge915 (.CLK_N(clknet_4_13_0_clk),
    .D(net707),
    .RESET_B(net738),
    .Q(net810));
 sky130_fd_sc_hd__dfrtp_2 merge916 (.CLK(clknet_4_8_0_clk),
    .D(net510),
    .RESET_B(net502),
    .Q(net811));
 sky130_fd_sc_hd__dfrtp_4 merge917 (.CLK(clknet_4_7_0_clk),
    .D(net726),
    .RESET_B(net747),
    .Q(net812));
 sky130_fd_sc_hd__dfrtp_4 merge918 (.CLK(clknet_4_15_0_clk),
    .D(net63),
    .RESET_B(net674),
    .Q(net813));
 sky130_fd_sc_hd__dfsbp_1 merge919 (.CLK(clknet_4_9_0_clk),
    .D(net714),
    .SET_B(net656),
    .Q(net1012),
    .Q_N(net814));
 sky130_fd_sc_hd__dfsbp_1 merge920 (.CLK(clknet_4_11_0_clk),
    .D(net764),
    .SET_B(net731),
    .Q(net815),
    .Q_N(net966));
 sky130_fd_sc_hd__dfstp_2 merge921 (.CLK(clknet_4_14_0_clk),
    .D(net685),
    .SET_B(net724),
    .Q(net816));
 sky130_fd_sc_hd__dfstp_4 merge922 (.CLK(clknet_4_0_0_clk),
    .D(net582),
    .SET_B(net673),
    .Q(net817));
 sky130_fd_sc_hd__dfstp_4 merge923 (.CLK(clknet_4_4_0_clk),
    .D(net325),
    .SET_B(net384),
    .Q(net818));
 sky130_fd_sc_hd__dlrbn_1 merge924 (.D(net736),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net737),
    .Q(net820),
    .Q_N(net819));
 sky130_fd_sc_hd__dlrbn_1 merge925 (.D(net783),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net782),
    .Q(net822),
    .Q_N(net821));
 sky130_fd_sc_hd__dlrbp_1 merge926 (.D(net398),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net499),
    .Q(net823),
    .Q_N(net1013));
 sky130_fd_sc_hd__dlrbp_1 merge927 (.D(net518),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net756),
    .Q(net825),
    .Q_N(net824));
 sky130_fd_sc_hd__dlrtn_1 merge928 (.D(net517),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net762),
    .Q(net963));
 sky130_fd_sc_hd__dlrtn_1 merge929 (.D(net414),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net405),
    .Q(net977));
 sky130_fd_sc_hd__dfxbp_1 s930 (.CLK(clknet_4_15_0_clk),
    .D(net40),
    .Q(net827),
    .Q_N(net826));
 sky130_fd_sc_hd__dfxbp_1 s931 (.CLK(clknet_4_15_0_clk),
    .D(net68),
    .Q(net983),
    .Q_N(net828));
 sky130_fd_sc_hd__dfxtp_2 s932 (.CLK(clknet_4_7_0_clk),
    .D(net116),
    .Q(net829));
 sky130_fd_sc_hd__dfxtp_1 s933 (.CLK(clknet_4_7_0_clk),
    .D(net134),
    .Q(net830));
 sky130_fd_sc_hd__dfxtp_1 s934 (.CLK(clknet_4_7_0_clk),
    .D(net137),
    .Q(net831));
 sky130_fd_sc_hd__dlclkp_1 s935 (.CLK(clknet_4_12_0_clk),
    .GATE(net155),
    .GCLK(net832));
 sky130_fd_sc_hd__dlclkp_2 s936 (.CLK(clknet_4_12_0_clk),
    .GATE(net156),
    .GCLK(net992));
 sky130_fd_sc_hd__dlclkp_4 s937 (.CLK(clknet_4_15_0_clk),
    .GATE(net188),
    .GCLK(net1002));
 sky130_fd_sc_hd__dlxbn_1 s938 (.D(net219),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net834),
    .Q_N(net833));
 sky130_fd_sc_hd__dlxbn_2 s939 (.D(net222),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net960),
    .Q_N(net835));
 sky130_fd_sc_hd__dlxbp_1 s940 (.D(net243),
    .GATE(clknet_4_4_0_clk),
    .Q(net837),
    .Q_N(net836));
 sky130_fd_sc_hd__dlxtn_2 s941 (.D(net250),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net838));
 sky130_fd_sc_hd__dlxtn_2 s942 (.D(net253),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net839));
 sky130_fd_sc_hd__dlxtn_4 s943 (.D(net282),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net840));
 sky130_fd_sc_hd__dlxtp_1 s944 (.D(net285),
    .GATE(clknet_4_12_0_clk),
    .Q(net841));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s945 (.D(net288),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net842));
 sky130_fd_sc_hd__dfxbp_2 s946 (.CLK(clknet_4_14_0_clk),
    .D(net295),
    .Q(net844),
    .Q_N(net843));
 sky130_fd_sc_hd__dfxbp_1 s947 (.CLK(clknet_4_14_0_clk),
    .D(net299),
    .Q(net846),
    .Q_N(net845));
 sky130_fd_sc_hd__dfxtp_1 s948 (.CLK(clknet_4_14_0_clk),
    .D(net305),
    .Q(net980));
 sky130_fd_sc_hd__dfxtp_4 s949 (.CLK(clknet_4_4_0_clk),
    .D(net323),
    .Q(net990));
 sky130_fd_sc_hd__dfxtp_2 s950 (.CLK(clknet_4_4_0_clk),
    .D(net327),
    .Q(net847));
 sky130_fd_sc_hd__dlclkp_1 s951 (.CLK(clknet_4_4_0_clk),
    .GATE(net328),
    .GCLK(net848));
 sky130_fd_sc_hd__dlclkp_2 s952 (.CLK(clknet_4_4_0_clk),
    .GATE(net340),
    .GCLK(net849));
 sky130_fd_sc_hd__dlclkp_4 s953 (.CLK(clknet_4_4_0_clk),
    .GATE(net343),
    .GCLK(net850));
 sky130_fd_sc_hd__dlxbn_1 s954 (.D(net345),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net852),
    .Q_N(net851));
 sky130_fd_sc_hd__dlxbn_1 s955 (.D(net346),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net854),
    .Q_N(net853));
 sky130_fd_sc_hd__dlxbp_1 s956 (.D(net348),
    .GATE(clknet_4_6_0_clk),
    .Q(net856),
    .Q_N(net855));
 sky130_fd_sc_hd__dlxtn_1 s957 (.D(net368),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net857));
 sky130_fd_sc_hd__dlxtn_4 s958 (.D(net369),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net981));
 sky130_fd_sc_hd__dlxtn_1 s959 (.D(net406),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net858));
 sky130_fd_sc_hd__dlxtp_1 s960 (.D(net408),
    .GATE(clknet_4_14_0_clk),
    .Q(net859));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s961 (.D(net412),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net860));
 sky130_fd_sc_hd__dfxbp_1 s962 (.CLK(clknet_4_1_0_clk),
    .D(net435),
    .Q(net862),
    .Q_N(net861));
 sky130_fd_sc_hd__dfxbp_1 s963 (.CLK(clknet_4_3_0_clk),
    .D(net472),
    .Q(net864),
    .Q_N(net863));
 sky130_fd_sc_hd__dfxtp_2 s964 (.CLK(clknet_4_3_0_clk),
    .D(net474),
    .Q(net865));
 sky130_fd_sc_hd__dfxtp_4 s965 (.CLK(clknet_4_3_0_clk),
    .D(net475),
    .Q(net866));
 sky130_fd_sc_hd__dfxtp_4 s966 (.CLK(clknet_4_3_0_clk),
    .D(net482),
    .Q(net867));
 sky130_fd_sc_hd__dlclkp_1 s967 (.CLK(clknet_4_3_0_clk),
    .GATE(net486),
    .GCLK(net868));
 sky130_fd_sc_hd__dlclkp_2 s968 (.CLK(clknet_4_3_0_clk),
    .GATE(net490),
    .GCLK(net869));
 sky130_fd_sc_hd__dlclkp_4 s969 (.CLK(clknet_4_3_0_clk),
    .GATE(net493),
    .GCLK(net969));
 sky130_fd_sc_hd__dlxbn_2 s970 (.D(net505),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net871),
    .Q_N(net870));
 sky130_fd_sc_hd__dlxbn_1 s971 (.D(net507),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net873),
    .Q_N(net872));
 sky130_fd_sc_hd__dlxbp_1 s972 (.D(net512),
    .GATE(clknet_4_10_0_clk),
    .Q(net875),
    .Q_N(net874));
 sky130_fd_sc_hd__dlxtn_1 s973 (.D(net524),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net973));
 sky130_fd_sc_hd__dlxtn_1 s974 (.D(net526),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net876));
 sky130_fd_sc_hd__dlxtn_1 s975 (.D(net529),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net877));
 sky130_fd_sc_hd__dlxtp_1 s976 (.D(net531),
    .GATE(clknet_4_10_0_clk),
    .Q(net878));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s977 (.D(net544),
    .SLEEP_B(clknet_4_0_0_clk),
    .Q(net879));
 sky130_fd_sc_hd__dfxbp_2 s978 (.CLK(clknet_4_2_0_clk),
    .D(net563),
    .Q(net881),
    .Q_N(net880));
 sky130_fd_sc_hd__dfxbp_2 s979 (.CLK(clknet_4_2_0_clk),
    .D(net571),
    .Q(net883),
    .Q_N(net882));
 sky130_fd_sc_hd__dfxtp_1 s980 (.CLK(clknet_4_2_0_clk),
    .D(net583),
    .Q(net884));
 sky130_fd_sc_hd__dfxtp_1 s981 (.CLK(clknet_4_2_0_clk),
    .D(net592),
    .Q(net885));
 sky130_fd_sc_hd__dfxtp_1 s982 (.CLK(clknet_4_2_0_clk),
    .D(net600),
    .Q(net886));
 sky130_fd_sc_hd__dlclkp_1 s983 (.CLK(clknet_4_8_0_clk),
    .GATE(net609),
    .GCLK(net887));
 sky130_fd_sc_hd__dlclkp_2 s984 (.CLK(clknet_4_2_0_clk),
    .GATE(net610),
    .GCLK(net888));
 sky130_fd_sc_hd__dlclkp_4 s985 (.CLK(clknet_4_8_0_clk),
    .GATE(net614),
    .GCLK(net889));
 sky130_fd_sc_hd__dlxbn_2 s986 (.D(net620),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net891),
    .Q_N(net890));
 sky130_fd_sc_hd__dlxbn_1 s987 (.D(net626),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net893),
    .Q_N(net892));
 sky130_fd_sc_hd__dlxbp_1 s988 (.D(net627),
    .GATE(clknet_4_8_0_clk),
    .Q(net895),
    .Q_N(net894));
 sky130_fd_sc_hd__dlxtn_2 s989 (.D(net635),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net896));
 sky130_fd_sc_hd__dlxtn_1 s990 (.D(net637),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net897));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in0),
    .X(net898));
 sky130_fd_sc_hd__buf_4 input2 (.A(in1),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(in10),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in12),
    .X(net902));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(in13),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net905));
 sky130_fd_sc_hd__buf_2 input9 (.A(in16),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in19),
    .X(net909));
 sky130_fd_sc_hd__buf_1 input13 (.A(in2),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net912));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(in23),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net916));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(in26),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net918));
 sky130_fd_sc_hd__buf_1 input22 (.A(in28),
    .X(net919));
 sky130_fd_sc_hd__buf_4 input23 (.A(in29),
    .X(net920));
 sky130_fd_sc_hd__buf_8 input24 (.A(in3),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_8 input26 (.A(in31),
    .X(net923));
 sky130_fd_sc_hd__buf_1 input27 (.A(in32),
    .X(net924));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(in34),
    .X(net926));
 sky130_fd_sc_hd__buf_4 input30 (.A(in35),
    .X(net927));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(in36),
    .X(net928));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(in38),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(in39),
    .X(net931));
 sky130_fd_sc_hd__buf_1 input35 (.A(in4),
    .X(net932));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net933));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in42),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net936));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net937));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net939));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net941));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net942));
 sky130_fd_sc_hd__buf_1 input46 (.A(in5),
    .X(net943));
 sky130_fd_sc_hd__buf_1 input47 (.A(in50),
    .X(net944));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(in52),
    .X(net946));
 sky130_fd_sc_hd__buf_1 input50 (.A(in53),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net948));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(in55),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(in56),
    .X(net950));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net951));
 sky130_fd_sc_hd__buf_4 input55 (.A(in58),
    .X(net952));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(in59),
    .X(net953));
 sky130_fd_sc_hd__buf_1 input57 (.A(in6),
    .X(net954));
 sky130_fd_sc_hd__buf_1 input58 (.A(in60),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(in61),
    .X(net956));
 sky130_fd_sc_hd__buf_2 input60 (.A(in7),
    .X(net957));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(in8),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(in9),
    .X(net959));
 sky130_fd_sc_hd__buf_2 output63 (.A(net960),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(clknet_1_1__leaf_net961),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net1058),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net963),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output67 (.A(net964),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output68 (.A(net965),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net966),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(clknet_1_0__leaf_net967),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net968),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(clknet_1_1__leaf_net969),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net970),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output74 (.A(net1020),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output75 (.A(net972),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output76 (.A(net973),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output77 (.A(net974),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output78 (.A(net975),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output79 (.A(net976),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output80 (.A(net977),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(clknet_1_0__leaf_net978),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output82 (.A(net979),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output83 (.A(net980),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output84 (.A(net981),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net982),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output86 (.A(net983),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output87 (.A(net984),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output88 (.A(net1018),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(clknet_1_1__leaf_net986),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output90 (.A(net987),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output91 (.A(net988),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output92 (.A(net989),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output93 (.A(net990),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net991),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(clknet_1_0__leaf_net992),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(clknet_1_1__leaf_net993),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output97 (.A(net994),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output98 (.A(net995),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output99 (.A(net996),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output100 (.A(net997),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(clknet_1_1__leaf_net998),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output102 (.A(net999),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net1000),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output104 (.A(net1001),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(clknet_1_1__leaf_net1002),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net1003),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output107 (.A(net1004),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output108 (.A(net1005),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output109 (.A(net1006),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output110 (.A(net1007),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(clknet_1_1__leaf_net1008),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output112 (.A(net1009),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(clknet_1_1__leaf_net1010),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output114 (.A(net1011),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output115 (.A(net1012),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output116 (.A(net1013),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(net982),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net1017),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net309),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_2 max_cap121 (.A(net985),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net1006),
    .X(net1019));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net971),
    .X(net1020));
 sky130_fd_sc_hd__buf_1 max_cap124 (.A(net211),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net5),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_2 wire126 (.A(net266),
    .X(net1023));
 sky130_fd_sc_hd__buf_2 wire127 (.A(net257),
    .X(net1024));
 sky130_fd_sc_hd__buf_1 max_cap128 (.A(net60),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net535),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net1028),
    .X(net1027));
 sky130_fd_sc_hd__buf_2 fanout131 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net457),
    .X(net1029));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(net333),
    .X(net1030));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net98),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_4 max_cap135 (.A(net860),
    .X(net1032));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(net319),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net1036),
    .X(net1035));
 sky130_fd_sc_hd__clkbuf_2 fanout139 (.A(net1039),
    .X(net1036));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net1039),
    .X(net1037));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net1039),
    .X(net1038));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net94),
    .X(net1039));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(net72),
    .X(net1040));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(net71),
    .X(net1041));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net58),
    .X(net1042));
 sky130_fd_sc_hd__buf_6 fanout146 (.A(net906),
    .X(net1043));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(net941),
    .X(net1044));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net924),
    .X(net1045));
 sky130_fd_sc_hd__inv_16 c192_1 (.A(clknet_1_0__leaf_net769),
    .Y(net1046));
 sky130_fd_sc_hd__clkinv_2 c214_3 (.A(net771),
    .Y(net1048));
 sky130_fd_sc_hd__clkinv_8 c79_5 (.A(net771),
    .Y(net1050));
 sky130_fd_sc_hd__clkinv_8 c79_6 (.A(net771),
    .Y(net1051));
 sky130_fd_sc_hd__clkinv_8 c79_7 (.A(net771),
    .Y(net1052));
 sky130_fd_sc_hd__inv_4 c85_9 (.A(net771),
    .Y(net1054));
 sky130_fd_sc_hd__inv_4 c85_10 (.A(net771),
    .Y(net1055));
 sky130_fd_sc_hd__clkinv_2 c352_14 (.A(net804),
    .Y(net1059));
 sky130_fd_sc_hd__clkinv_2 c352_15 (.A(net804),
    .Y(net1060));
 sky130_fd_sc_hd__clkinv_2 c352_16 (.A(net804),
    .Y(net1061));
 sky130_fd_sc_hd__clkinv_2 c352_17 (.A(net804),
    .Y(net1062));
 sky130_fd_sc_hd__clkinv_2 c352_18 (.A(net804),
    .Y(net1063));
 sky130_fd_sc_hd__clkinv_2 c352_19 (.A(net804),
    .Y(net1064));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net889 (.A(net889),
    .X(clknet_0_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net889 (.A(clknet_0_net889),
    .X(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net889 (.A(clknet_0_net889),
    .X(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net888 (.A(net888),
    .X(clknet_0_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net888 (.A(clknet_0_net888),
    .X(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net888 (.A(clknet_0_net888),
    .X(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net770 (.A(net770),
    .X(clknet_0_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net770 (.A(clknet_0_net770),
    .X(clknet_1_0__leaf_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net770 (.A(clknet_0_net770),
    .X(clknet_1_1__leaf_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net617 (.A(net617),
    .X(clknet_0_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_0__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_1__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net887 (.A(net887),
    .X(clknet_0_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net612 (.A(net612),
    .X(clknet_0_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net612 (.A(clknet_0_net612),
    .X(clknet_1_0__leaf_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net612 (.A(clknet_0_net612),
    .X(clknet_1_1__leaf_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net616 (.A(net616),
    .X(clknet_0_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_0__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_1__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net969 (.A(net969),
    .X(clknet_0_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_0__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_1__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net869 (.A(net869),
    .X(clknet_0_net869));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net869 (.A(clknet_0_net869),
    .X(clknet_1_0__leaf_net869));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net869 (.A(clknet_0_net869),
    .X(clknet_1_1__leaf_net869));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net504 (.A(net504),
    .X(clknet_0_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_0__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_1__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net868 (.A(net868),
    .X(clknet_0_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_1__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net850 (.A(net850),
    .X(clknet_0_net850));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net850 (.A(clknet_0_net850),
    .X(clknet_1_0__leaf_net850));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net850 (.A(clknet_0_net850),
    .X(clknet_1_1__leaf_net850));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net356 (.A(net356),
    .X(clknet_0_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_0__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_1__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net351 (.A(net351),
    .X(clknet_0_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_0__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_1__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net978 (.A(net978),
    .X(clknet_0_net978));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net978 (.A(clknet_0_net978),
    .X(clknet_1_0__leaf_net978));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net978 (.A(clknet_0_net978),
    .X(clknet_1_1__leaf_net978));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net849 (.A(net849),
    .X(clknet_0_net849));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net849 (.A(clknet_0_net849),
    .X(clknet_1_0__leaf_net849));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net849 (.A(clknet_0_net849),
    .X(clknet_1_1__leaf_net849));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net342 (.A(net342),
    .X(clknet_0_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net848 (.A(net848),
    .X(clknet_0_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net848 (.A(clknet_0_net848),
    .X(clknet_1_0__leaf_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net848 (.A(clknet_0_net848),
    .X(clknet_1_1__leaf_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net541 (.A(net541),
    .X(clknet_0_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_0__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_1__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net546 (.A(net546),
    .X(clknet_0_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net546 (.A(clknet_0_net546),
    .X(clknet_1_0__leaf_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net546 (.A(clknet_0_net546),
    .X(clknet_1_1__leaf_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net418 (.A(net418),
    .X(clknet_0_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net418 (.A(clknet_0_net418),
    .X(clknet_1_0__leaf_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net418 (.A(clknet_0_net418),
    .X(clknet_1_1__leaf_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net432 (.A(net432),
    .X(clknet_0_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net432 (.A(clknet_0_net432),
    .X(clknet_1_0__leaf_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net432 (.A(clknet_0_net432),
    .X(clknet_1_1__leaf_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net536 (.A(net536),
    .X(clknet_0_net536));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net536 (.A(clknet_0_net536),
    .X(clknet_1_0__leaf_net536));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net536 (.A(clknet_0_net536),
    .X(clknet_1_1__leaf_net536));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net438 (.A(net438),
    .X(clknet_0_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_0__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_1__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net429 (.A(net429),
    .X(clknet_0_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_1__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net485 (.A(net485),
    .X(clknet_0_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_0__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_1__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net464 (.A(net464),
    .X(clknet_0_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net427 (.A(net427),
    .X(clknet_0_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_1__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net445 (.A(net445),
    .X(clknet_0_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_0__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_1__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net967 (.A(net967),
    .X(clknet_0_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net967 (.A(clknet_0_net967),
    .X(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net967 (.A(clknet_0_net967),
    .X(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net503 (.A(net503),
    .X(clknet_0_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_1__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net425 (.A(net425),
    .X(clknet_0_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_0__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_1__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net430 (.A(net430),
    .X(clknet_0_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_0__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_1__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net417 (.A(net417),
    .X(clknet_0_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net417 (.A(clknet_0_net417),
    .X(clknet_1_0__leaf_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net417 (.A(clknet_0_net417),
    .X(clknet_1_1__leaf_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1002 (.A(net1002),
    .X(clknet_0_net1002));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1002 (.A(clknet_0_net1002),
    .X(clknet_1_0__leaf_net1002));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1002 (.A(clknet_0_net1002),
    .X(clknet_1_1__leaf_net1002));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net190 (.A(net190),
    .X(clknet_0_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net190 (.A(clknet_0_net190),
    .X(clknet_1_0__leaf_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net190 (.A(clknet_0_net190),
    .X(clknet_1_1__leaf_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net993 (.A(net993),
    .X(clknet_0_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net993 (.A(clknet_0_net993),
    .X(clknet_1_0__leaf_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net993 (.A(clknet_0_net993),
    .X(clknet_1_1__leaf_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net992 (.A(net992),
    .X(clknet_0_net992));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net992 (.A(clknet_0_net992),
    .X(clknet_1_0__leaf_net992));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net992 (.A(clknet_0_net992),
    .X(clknet_1_1__leaf_net992));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net832 (.A(net832),
    .X(clknet_0_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net832 (.A(clknet_0_net832),
    .X(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net832 (.A(clknet_0_net832),
    .X(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net371 (.A(net371),
    .X(clknet_0_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_0__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_1__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net374 (.A(net374),
    .X(clknet_0_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net374 (.A(clknet_0_net374),
    .X(clknet_1_0__leaf_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net374 (.A(clknet_0_net374),
    .X(clknet_1_1__leaf_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net986 (.A(net986),
    .X(clknet_0_net986));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net986 (.A(clknet_0_net986),
    .X(clknet_1_0__leaf_net986));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net986 (.A(clknet_0_net986),
    .X(clknet_1_1__leaf_net986));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net36 (.A(net36),
    .X(clknet_0_net36));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net36 (.A(clknet_0_net36),
    .X(clknet_1_0__leaf_net36));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net36 (.A(clknet_0_net36),
    .X(clknet_1_1__leaf_net36));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net38 (.A(net38),
    .X(clknet_0_net38));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net38 (.A(clknet_0_net38),
    .X(clknet_1_0__leaf_net38));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net38 (.A(clknet_0_net38),
    .X(clknet_1_1__leaf_net38));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net35 (.A(net35),
    .X(clknet_0_net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net35 (.A(clknet_0_net35),
    .X(clknet_1_0__leaf_net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net35 (.A(clknet_0_net35),
    .X(clknet_1_1__leaf_net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net39 (.A(net39),
    .X(clknet_0_net39));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net39 (.A(clknet_0_net39),
    .X(clknet_1_0__leaf_net39));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net39 (.A(clknet_0_net39),
    .X(clknet_1_1__leaf_net39));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net998 (.A(net998),
    .X(clknet_0_net998));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net998 (.A(clknet_0_net998),
    .X(clknet_1_0__leaf_net998));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net998 (.A(clknet_0_net998),
    .X(clknet_1_1__leaf_net998));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net304 (.A(net304),
    .X(clknet_0_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net304 (.A(clknet_0_net304),
    .X(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net304 (.A(clknet_0_net304),
    .X(clknet_1_1__leaf_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net516 (.A(net516),
    .X(clknet_0_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_0__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_1__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net172 (.A(net172),
    .X(clknet_0_net172));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net172 (.A(clknet_0_net172),
    .X(clknet_1_0__leaf_net172));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net172 (.A(clknet_0_net172),
    .X(clknet_1_1__leaf_net172));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net175 (.A(net175),
    .X(clknet_0_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_0__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_1__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net176 (.A(net176),
    .X(clknet_0_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net176 (.A(clknet_0_net176),
    .X(clknet_1_0__leaf_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net176 (.A(clknet_0_net176),
    .X(clknet_1_1__leaf_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net168 (.A(net168),
    .X(clknet_0_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_0__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_1__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net961 (.A(net961),
    .X(clknet_0_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net961 (.A(clknet_0_net961),
    .X(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net961 (.A(clknet_0_net961),
    .X(clknet_1_1__leaf_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net167 (.A(net167),
    .X(clknet_0_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_0__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_1__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net24 (.A(net24),
    .X(clknet_0_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net24 (.A(clknet_0_net24),
    .X(clknet_1_0__leaf_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net24 (.A(clknet_0_net24),
    .X(clknet_1_1__leaf_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net25 (.A(net25),
    .X(clknet_0_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net25 (.A(clknet_0_net25),
    .X(clknet_1_0__leaf_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net25 (.A(clknet_0_net25),
    .X(clknet_1_1__leaf_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net54 (.A(net54),
    .X(clknet_0_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net54 (.A(clknet_0_net54),
    .X(clknet_1_0__leaf_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net54 (.A(clknet_0_net54),
    .X(clknet_1_1__leaf_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net19 (.A(net19),
    .X(clknet_0_net19));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net19 (.A(clknet_0_net19),
    .X(clknet_1_0__leaf_net19));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net19 (.A(clknet_0_net19),
    .X(clknet_1_1__leaf_net19));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1010 (.A(net1010),
    .X(clknet_0_net1010));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1010 (.A(clknet_0_net1010),
    .X(clknet_1_0__leaf_net1010));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1010 (.A(clknet_0_net1010),
    .X(clknet_1_1__leaf_net1010));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net22 (.A(net22),
    .X(clknet_0_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net22 (.A(clknet_0_net22),
    .X(clknet_1_0__leaf_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net22 (.A(clknet_0_net22),
    .X(clknet_1_1__leaf_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net140 (.A(net140),
    .X(clknet_0_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_0__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net29 (.A(net29),
    .X(clknet_0_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net29 (.A(clknet_0_net29),
    .X(clknet_1_0__leaf_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net29 (.A(clknet_0_net29),
    .X(clknet_1_1__leaf_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net34 (.A(net34),
    .X(clknet_0_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net34 (.A(clknet_0_net34),
    .X(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net34 (.A(clknet_0_net34),
    .X(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net30 (.A(net30),
    .X(clknet_0_net30));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net30 (.A(clknet_0_net30),
    .X(clknet_1_0__leaf_net30));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net30 (.A(clknet_0_net30),
    .X(clknet_1_1__leaf_net30));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net769 (.A(net769),
    .X(clknet_0_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_1__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net12 (.A(net12),
    .X(clknet_0_net12));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net12 (.A(clknet_0_net12),
    .X(clknet_1_0__leaf_net12));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net12 (.A(clknet_0_net12),
    .X(clknet_1_1__leaf_net12));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net16 (.A(net16),
    .X(clknet_0_net16));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net16 (.A(clknet_0_net16),
    .X(clknet_1_0__leaf_net16));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net16 (.A(clknet_0_net16),
    .X(clknet_1_1__leaf_net16));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net303 (.A(net303),
    .X(clknet_0_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_0__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_1__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net169 (.A(net169),
    .X(clknet_0_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net157 (.A(net157),
    .X(clknet_0_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_1__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1008 (.A(net1008),
    .X(clknet_0_net1008));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1008 (.A(clknet_0_net1008),
    .X(clknet_1_0__leaf_net1008));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1008 (.A(clknet_0_net1008),
    .X(clknet_1_1__leaf_net1008));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net130 (.A(net130),
    .X(clknet_0_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_1__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net111 (.A(net111),
    .X(clknet_0_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_0__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_1__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net110 (.A(net110),
    .X(clknet_0_net110));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net110 (.A(clknet_0_net110),
    .X(clknet_1_0__leaf_net110));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net110 (.A(clknet_0_net110),
    .X(clknet_1_1__leaf_net110));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net1098),
    .X(net17));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net17),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net17),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net338),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1098),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net338),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net746),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net729),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net847),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net538),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net396),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net545),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net48),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net173),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net794),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net833),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net865),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net41),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net846),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net761),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net772),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net161),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net980),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net837),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net312),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net89),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net215),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net61),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net153),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net979),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net976),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net806),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net786),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net556),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net125),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net886),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net255),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net884),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net113),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net828),
    .X(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_A3 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_A0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_C1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_X (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_C (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_C (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A3 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SCD (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_C1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_Y (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_C (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_Y (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_C1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_SCD (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_Y (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_A3 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_C (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold29_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_Y (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_Y (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_S0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_X (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_Y (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_RESET_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_C1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_D (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A3 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_SCE (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_S1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_SCE (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_Y (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_C_N (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Y (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_C1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_Y (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A_N (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_S0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A_N (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_SCE (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Y (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold27_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_SCD (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_S0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_Q_N (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_Q (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B_N (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Y (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_S1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_SCE (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_SCD (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCE (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_Y (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_C_N (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_DE (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_X (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_C_N (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A_N (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_DE (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_Q (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A3 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_Y (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_SCE (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_Y (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_Y (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_C1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_Q_N (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_Q (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_S1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SCD (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Y (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_D (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_D (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B_N (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_DE (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_Y (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_Q (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Q (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_B1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B2 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_RESET_B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A3 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B_N (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_DE (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_Y (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_Q_N (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_B2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_RESET_B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_Y (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCE (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SCE (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_X (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net374_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_X (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge923_SET_B (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_X (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_RESET_B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_B2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_Y (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_Y (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_SCE (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_Q_N (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_C (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_Q (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SCD (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_C (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_Y (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_C (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_Q_N (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCD (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_C (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_B2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_SCD (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_X (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A3 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_Q_N (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_Q (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_S1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_A3 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_Y (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_X (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_S1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_SET_B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_SCD (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S0 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_RESET_B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_X (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SCD (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_X (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net546_A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_Y (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_B2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_SCD (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_X (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_B1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SCE (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_B1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_Q (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_Q (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_B2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_Y (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge896_SET_B (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_X (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge921_D (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_Y (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_D (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_Y (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_Q (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_C1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold20_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_Q (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_Q (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_C1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_10_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_9_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_8_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_7_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_6_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_5_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_4_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_3_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_2_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_GCLK (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_Q (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_Q (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_Q (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_C1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_SCD (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCD (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_SCE (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Y (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge895_Q (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge905_Q (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_B2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge906_Q (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_B2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_Y (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_Y (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge909_Q (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_19_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_18_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_17_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_16_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_15_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_14_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_13_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge911_GCLK (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_SCE (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge915_Q (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_SCE (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge917_Q (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_C1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SET_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_C (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_C1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_C_N (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge918_Q (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge921_Q (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge923_Q (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_C1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_C (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_C1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_Q (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A_N (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_C1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_Y (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_Q_N (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_Q (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_C (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_C (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_Q (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_C1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_C_N (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_C1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_Q (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A_N (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_SCD (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_s962_Q (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_C1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_s965_Q (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_B2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_B2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_Q (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_B1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_s970_Q (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_s971_Q (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_s978_Q_N (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_B2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold38_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_s980_Q (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_Q (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A3 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_Y (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_Y (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCD (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_B2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_C (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A_N (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_A0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B_N (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_C_N (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_C1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A3 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A3 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_S1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B_N (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_D (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B_N (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A_N (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_C1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_C1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_SCE (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_C1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_SCD (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_SCD (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A_N (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_D (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A3 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_SCE (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_B1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_C1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_D (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_Q (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge928_Q (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_Q (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_SCE (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_Y (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_Y (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCD (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_Q (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_Q (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge929_Q (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_Q (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_B1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_Y (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap121_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_SCE (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_SCD (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_Y (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_Q (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_C1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_Y (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_D (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_Y (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_Q (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net992_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_GCLK (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_Y (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_Y (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_SCD (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_RESET_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_Q (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_C1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_SCD (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_C1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_C_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_B1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_C1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_Y (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_Y (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net1008_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_Y (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_Q (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge919_Q (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_C1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge926_Q_N (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_C_N (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_C1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_S0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_SCD (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_SCD (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_C1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_S1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap121_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_SCE (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_SET_B (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_B2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_RESET_B (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_SCE (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_D (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SCD (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire127_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCD (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_C1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCE (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_SET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_SET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_C1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_C1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_C1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_SCE (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SCD (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_SCE (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_C1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_S1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_SCD (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap135_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A_N (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_SCD (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_B1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_B2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_C (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SCE (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_C (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B_N (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_S0 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SCE (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_C (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCE (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_C (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_C (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_C (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A_N (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_RESET_B (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_S1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_C (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B_N (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_B1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_C1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S0 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SCD (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge900_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge922_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s977_SLEEP_B (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge913_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s954_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s962_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge902_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s978_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s979_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s980_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s981_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s982_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s984_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge906_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge907_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge908_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge910_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s965_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s968_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s969_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge904_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge923_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge897_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s956_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge917_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge924_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge896_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge916_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge925_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s970_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s971_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s983_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s985_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s986_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s987_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s988_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge905_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge914_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge919_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge928_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge892_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge920_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge926_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge929_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s974_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge895_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge901_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge899_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge915_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge911_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge921_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_SLEEP_B (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_SLEEP_B (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge891_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge898_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge918_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_C1 (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net868_X (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(clknet_1_0__leaf_net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(clknet_1_0__leaf_net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net978_X (.DIODE(clknet_1_0__leaf_net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S1 (.DIODE(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SCE (.DIODE(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_A2 (.DIODE(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net429_X (.DIODE(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A1 (.DIODE(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net464_X (.DIODE(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net464_X (.DIODE(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_12_A (.DIODE(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net967_X (.DIODE(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_B (.DIODE(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_11_A (.DIODE(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net967_X (.DIODE(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(clknet_1_0__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(clknet_1_0__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(clknet_1_0__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(clknet_1_0__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net992_X (.DIODE(clknet_1_0__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(clknet_1_1__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(clknet_1_1__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(clknet_1_1__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(clknet_1_1__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net992_X (.DIODE(clknet_1_1__leaf_net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_RESET_B (.DIODE(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net961_X (.DIODE(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_C1 (.DIODE(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCD (.DIODE(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_C1 (.DIODE(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net34_X (.DIODE(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_RESET_B (.DIODE(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A1 (.DIODE(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net34_X (.DIODE(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net162_X (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_RESET_B (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_X (.DIODE(net1075));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net338),
    .X(net1098));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
