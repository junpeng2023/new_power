module netlist_0 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input in52,
	input in53,
	input in54,
	input in55,
	input in56,
	input in57,
	input in58,
	input in59,
	input in60,
	input in61,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51,
	output out52,
	output out53,
	output out54,
	output out55,
	output out56,
	output out57,
	output out58,
	output out59,
	output out60,
	output out61
);


wire clk;
wire out3;
wire net825;
wire net823;
wire net822;
wire net821;
wire net820;
wire net819;
wire net818;
wire net817;
wire net816;
wire net815;
wire net814;
wire net813;
wire net812;
wire net811;
wire net810;
wire net807;
wire net805;
wire net804;
wire net802;
wire net801;
wire net800;
wire net795;
wire out2;
wire net793;
wire net792;
wire net791;
wire net789;
wire out20;
wire net787;
wire net786;
wire net785;
wire net784;
wire out17;
wire net808;
wire net781;
wire net780;
wire net777;
wire net776;
wire out1;
wire net775;
wire net774;
wire net773;
wire net772;
wire net771;
wire net770;
wire net769;
wire net766;
wire net765;
wire net764;
wire out53;
wire net763;
wire net762;
wire out19;
wire out30;
wire net759;
wire net755;
wire net754;
wire out35;
wire net753;
wire net752;
wire net751;
wire net750;
wire out11;
wire net748;
wire net790;
wire net747;
wire net745;
wire net744;
wire net743;
wire net741;
wire net740;
wire net739;
wire net738;
wire net735;
wire net732;
wire out42;
wire net731;
wire net730;
wire out13;
wire net729;
wire net728;
wire net726;
wire net725;
wire net724;
wire net722;
wire net720;
wire net719;
wire net717;
wire net716;
wire net715;
wire net714;
wire net712;
wire net711;
wire net708;
wire net706;
wire net705;
wire net704;
wire out16;
wire net703;
wire net701;
wire net699;
wire net779;
wire net698;
wire out49;
wire net692;
wire net690;
wire net299;
wire net688;
wire net686;
wire net684;
wire net683;
wire out57;
wire net503;
wire net679;
wire net671;
wire net669;
wire net668;
wire net370;
wire net667;
wire net664;
wire net694;
wire net659;
wire in6;
wire net656;
wire net652;
wire net622;
wire net651;
wire net304;
wire net645;
wire net641;
wire net637;
wire net632;
wire net665;
wire net631;
wire net629;
wire net74;
wire net628;
wire net3;
wire net627;
wire net447;
wire net626;
wire net624;
wire net506;
wire net623;
wire net620;
wire in49;
wire net619;
wire net798;
wire net46;
wire net615;
wire net347;
wire net100;
wire net288;
wire net614;
wire net165;
wire net613;
wire net20;
wire net612;
wire net638;
wire net428;
wire net610;
wire out25;
wire net608;
wire net1;
wire net424;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire net782;
wire net601;
wire net596;
wire net592;
wire net588;
wire net587;
wire in4;
wire net583;
wire net707;
wire net582;
wire net158;
wire net584;
wire net581;
wire net336;
wire net579;
wire net577;
wire net576;
wire net570;
wire net209;
wire net569;
wire in41;
wire net567;
wire net696;
wire net794;
wire in30;
wire net566;
wire net565;
wire net39;
wire net562;
wire net559;
wire net556;
wire net647;
wire net555;
wire net159;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire in55;
wire net550;
wire net710;
wire net544;
wire net539;
wire net534;
wire net532;
wire net271;
wire net530;
wire net617;
wire net306;
wire net537;
wire net369;
wire net528;
wire net525;
wire net523;
wire net520;
wire net519;
wire net516;
wire net672;
wire net514;
wire net512;
wire net78;
wire net508;
wire net721;
wire net504;
wire net224;
wire net573;
wire net499;
wire net674;
wire net496;
wire net495;
wire net494;
wire net179;
wire in39;
wire net453;
wire net493;
wire net788;
wire net472;
wire net492;
wire net479;
wire net491;
wire net295;
wire net490;
wire net489;
wire net487;
wire net486;
wire net478;
wire net474;
wire net473;
wire net468;
wire net540;
wire net202;
wire net465;
wire out7;
wire net462;
wire net469;
wire net471;
wire net461;
wire net546;
wire net749;
wire net460;
wire net454;
wire net44;
wire net117;
wire net689;
wire net648;
wire net452;
wire net449;
wire net448;
wire net498;
wire net700;
wire net446;
wire net680;
wire net88;
wire net691;
wire net444;
wire in59;
wire net110;
wire net442;
wire net609;
wire net440;
wire net128;
wire net439;
wire out23;
wire out21;
wire net147;
wire net438;
wire net797;
wire net433;
wire net432;
wire out41;
wire net419;
wire net431;
wire net430;
wire net618;
wire net429;
wire net427;
wire net809;
wire net426;
wire net673;
wire net425;
wire net423;
wire net183;
wire net531;
wire net421;
wire net52;
wire net170;
wire net420;
wire net450;
wire net418;
wire net415;
wire net414;
wire net276;
wire net413;
wire net252;
wire net330;
wire net412;
wire net411;
wire net517;
wire net677;
wire net410;
wire net409;
wire net685;
wire net407;
wire net406;
wire net662;
wire net405;
wire net607;
wire net526;
wire net404;
wire net29;
wire net403;
wire net383;
wire net663;
wire net402;
wire net106;
wire net572;
wire net401;
wire net399;
wire net398;
wire net476;
wire net396;
wire net172;
wire net395;
wire net391;
wire net693;
wire net443;
wire net557;
wire net345;
wire net527;
wire net488;
wire net390;
wire out5;
wire net646;
wire net389;
wire net513;
wire net501;
wire out14;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net184;
wire net131;
wire net380;
wire net379;
wire net260;
wire net616;
wire net378;
wire net543;
wire net38;
wire net377;
wire net376;
wire net625;
wire net373;
wire net598;
wire net374;
wire net676;
wire net372;
wire net371;
wire out54;
wire net368;
wire net367;
wire net366;
wire net365;
wire net364;
wire net363;
wire net360;
wire net397;
wire net357;
wire net356;
wire net510;
wire net355;
wire net521;
wire net353;
wire net590;
wire net507;
wire net351;
wire net746;
wire net350;
wire net547;
wire net511;
wire net451;
wire net13;
wire net343;
wire net89;
wire net666;
wire net340;
wire net339;
wire net337;
wire net458;
wire net538;
wire net244;
wire net334;
wire net333;
wire net332;
wire net331;
wire out32;
wire net328;
wire net327;
wire net119;
wire net325;
wire net324;
wire out56;
wire net321;
wire out58;
wire net535;
wire net320;
wire out46;
wire net542;
wire net139;
wire net318;
wire net505;
wire net199;
wire out27;
wire net294;
wire net319;
wire net312;
wire net636;
wire net518;
wire in37;
wire net311;
wire net309;
wire net742;
wire net308;
wire net417;
wire out8;
wire net302;
wire net298;
wire net296;
wire in24;
wire net358;
wire net127;
wire net180;
wire net310;
wire net697;
wire net293;
wire net305;
wire net594;
wire out39;
wire net292;
wire net500;
wire net445;
wire net303;
wire net291;
wire net201;
wire net422;
wire net289;
wire net595;
wire net384;
wire net482;
wire in25;
wire net589;
wire net278;
wire net761;
wire net274;
wire net643;
wire net273;
wire net142;
wire out10;
wire net272;
wire net114;
wire net270;
wire in17;
wire net267;
wire net644;
wire net266;
wire out38;
wire net459;
wire net463;
wire net0;
wire net297;
wire net408;
wire net475;
wire net280;
wire net102;
wire net799;
wire net151;
wire net275;
wire net264;
wire net657;
wire net591;
wire net196;
wire net262;
wire net217;
wire net261;
wire net21;
wire net257;
wire net62;
wire net109;
wire net254;
wire net203;
wire net253;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire net767;
wire net111;
wire net124;
wire net242;
wire in26;
wire net661;
wire net194;
wire net241;
wire net238;
wire net234;
wire net232;
wire out12;
wire net226;
wire net568;
wire net375;
wire net223;
wire net524;
wire net575;
wire net382;
wire net548;
wire net259;
wire out9;
wire net315;
wire net335;
wire net222;
wire in29;
wire net240;
wire net416;
wire net41;
wire net104;
wire net8;
wire out33;
wire net31;
wire net219;
wire net578;
wire net210;
wire net326;
wire net213;
wire net208;
wire net188;
wire net207;
wire net649;
wire net205;
wire net678;
wire net633;
wire net122;
wire net197;
wire net483;
wire net193;
wire net192;
wire net737;
wire net190;
wire net630;
wire in20;
wire net189;
wire net246;
wire net783;
wire net186;
wire net660;
wire net359;
wire out28;
wire net152;
wire net126;
wire net113;
wire net284;
wire net655;
wire net563;
wire net464;
wire net549;
wire net182;
wire net258;
wire net176;
wire net580;
wire net133;
wire net175;
wire net80;
wire net173;
wire out52;
wire net195;
wire net381;
wire net218;
wire net300;
wire net169;
wire net485;
wire net344;
wire net168;
wire net153;
wire net286;
wire net167;
wire net509;
wire net58;
wire net221;
wire net166;
wire net269;
wire net97;
wire net434;
wire net204;
wire net200;
wire net621;
wire net162;
wire out60;
wire net497;
wire out45;
wire net161;
wire net285;
wire net160;
wire net149;
wire net695;
wire net148;
wire net178;
wire net239;
wire net144;
wire out31;
wire net316;
wire net322;
wire net758;
wire net143;
wire out37;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net806;
wire net561;
wire out29;
wire net137;
wire net136;
wire net456;
wire net135;
wire net255;
wire net157;
wire net177;
wire out48;
wire net134;
wire net150;
wire net441;
wire out15;
wire net130;
wire in12;
wire net103;
wire out18;
wire net481;
wire net120;
wire net455;
wire net65;
wire net129;
wire net392;
wire out0;
wire net164;
wire net687;
wire net642;
wire net268;
wire in7;
wire net756;
wire net400;
wire net82;
wire net2;
wire net123;
wire net282;
wire net71;
wire net229;
wire in43;
wire net108;
wire net107;
wire out26;
wire net99;
wire net348;
wire net341;
wire in52;
wire net96;
wire net225;
wire net250;
wire net466;
wire net118;
wire net94;
wire net90;
wire net803;
wire net174;
wire net277;
wire net639;
wire net81;
wire out22;
wire net230;
wire in10;
wire net156;
wire net361;
wire net115;
wire net670;
wire in18;
wire net27;
wire net34;
wire net585;
wire net79;
wire net75;
wire net231;
wire net349;
wire net329;
wire net212;
wire net653;
wire in5;
wire net14;
wire net77;
wire net600;
wire net236;
wire net76;
wire in42;
wire net354;
wire in38;
wire net736;
wire net198;
wire net467;
wire net101;
wire net9;
wire net571;
wire net73;
wire net116;
wire net69;
wire net67;
wire in31;
wire net98;
wire net522;
wire net436;
wire net541;
wire net323;
wire net15;
wire net279;
wire net64;
wire net63;
wire net681;
wire net61;
wire net60;
wire net682;
wire net237;
wire net59;
wire net248;
wire net477;
wire net564;
wire net154;
wire net84;
wire in46;
wire net85;
wire net72;
wire net228;
wire net675;
wire net56;
wire net55;
wire net214;
wire net53;
wire in48;
wire net640;
wire net50;
wire net597;
wire out55;
wire net185;
wire net155;
wire net338;
wire net599;
wire net112;
wire net650;
wire net560;
wire net45;
wire net502;
wire net235;
wire net49;
wire in50;
wire net215;
wire net484;
wire in8;
wire net346;
wire net4;
wire net43;
wire net187;
wire in13;
wire net586;
wire net533;
wire net796;
wire net32;
wire net125;
wire net19;
wire in15;
wire net727;
wire net163;
wire in19;
wire net702;
wire net70;
wire net48;
wire net28;
wire net92;
wire net713;
wire net25;
wire net30;
wire in0;
wire net709;
wire net24;
wire out47;
wire net290;
wire net227;
wire net470;
wire in33;
wire net33;
wire net824;
wire net233;
wire net121;
wire net40;
wire in60;
wire net435;
wire out34;
wire net18;
wire net301;
wire net760;
wire net23;
wire net26;
wire net16;
wire net558;
wire in1;
wire net265;
wire net778;
wire net22;
wire net263;
wire net457;
wire out50;
wire net6;
wire net5;
wire net206;
wire in58;
wire net342;
wire net17;
wire in61;
wire net757;
wire in56;
wire net733;
wire net171;
wire in23;
wire in51;
wire net317;
wire out4;
wire net42;
wire net91;
wire in57;
wire net281;
wire net54;
wire net313;
wire in54;
wire out43;
wire in53;
wire net138;
wire net145;
wire net211;
wire net132;
wire out24;
wire in35;
wire in34;
wire net593;
wire in45;
wire net393;
wire net256;
wire net87;
wire net181;
wire net7;
wire net574;
wire net216;
wire out59;
wire in28;
wire in44;
wire in32;
wire net47;
wire net12;
wire in27;
wire in9;
wire net654;
wire net723;
wire net611;
wire net515;
wire net362;
wire in16;
wire net191;
wire net35;
wire net220;
wire in22;
wire net68;
wire in14;
wire net529;
wire in21;
wire net57;
wire net480;
wire net86;
wire net93;
wire in47;
wire in2;
wire net718;
wire net658;
wire net105;
wire in11;
wire net51;
wire out44;
wire net437;
wire in36;
wire net536;
wire net37;
wire net36;
wire net95;
wire net146;
wire net394;
wire in3;
wire net314;
wire net734;
wire net251;
wire net768;
wire net11;
wire net352;
wire net307;
sky130_fd_sc_hd__mux4_2 c62(
.A0(in50),
.A1(in58),
.A2(in38),
.A3(in53),
.S0(in26),
.S1(in56),
.X(net0)
);

sky130_fd_sc_hd__mux4_1 c63(
.A0(in51),
.A1(in53),
.A2(in50),
.A3(net3),
.S0(in26),
.S1(in10),
.X(net1)
);

sky130_fd_sc_hd__mux4_1 c64(
.A0(in42),
.A1(in54),
.A2(in44),
.A3(in1),
.S0(in58),
.S1(in50),
.X(net2)
);

sky130_fd_sc_hd__mux4_1 c65(
.A0(in10),
.A1(in12),
.A2(in26),
.A3(in3),
.S0(in38),
.S1(in42),
.X(net3)
);

sky130_fd_sc_hd__nor2b_2 c66(
.A(in1),
.B_N(in46),
.Y(net4)
);

sky130_fd_sc_hd__and2b_2 c67(
.A_N(net4),
.B(in24),
.X(net5)
);

sky130_fd_sc_hd__or2_1 c68(
.A(in24),
.B(in45),
.X(net6)
);

sky130_fd_sc_hd__nor2_4 c69(
.A(in61),
.B(in38),
.Y(net7)
);

sky130_fd_sc_hd__nor2b_2 c70(
.A(in43),
.B_N(net1),
.Y(net8)
);

sky130_fd_sc_hd__a41o_4 c71(
.A1(in19),
.A2(in45),
.A3(net4),
.A4(in43),
.B1(in42),
.X(net9)
);

sky130_fd_sc_hd__nor2_4 c72(
.A(in20),
.B(in38),
.Y(net10)
);

sky130_fd_sc_hd__and2b_1 c73(
.A_N(net5),
.B(net10),
.X(net11)
);

sky130_fd_sc_hd__mux2_2 c74(
.A0(net10),
.A1(net8),
.S(in59),
.X(net12)
);

sky130_fd_sc_hd__nand2b_1 c75(
.A_N(in58),
.B(net7),
.Y(net13)
);

sky130_fd_sc_hd__or2_2 c76(
.A(net9),
.B(net11),
.X(net14)
);

sky130_fd_sc_hd__mux4_4 c77(
.A0(net6),
.A1(net4),
.A2(in36),
.A3(net11),
.S0(net8),
.S1(in46),
.X(net15)
);

sky130_fd_sc_hd__and2b_1 c78(
.A_N(net12),
.B(net15),
.X(net16)
);

sky130_fd_sc_hd__a31oi_4 c79(
.A1(net14),
.A2(net6),
.A3(net15),
.B1(net7),
.Y(net17)
);

sky130_fd_sc_hd__a31oi_2 c80(
.A1(net15),
.A2(net10),
.A3(in28),
.B1(in59),
.Y(net18)
);

sky130_fd_sc_hd__nor2_1 c81(
.A(in16),
.B(net2),
.Y(net19)
);

sky130_fd_sc_hd__a31o_2 c82(
.A1(in8),
.A2(net18),
.A3(in59),
.B1(net5),
.X(net20)
);

sky130_fd_sc_hd__mux4_1 c83(
.A0(net16),
.A1(net19),
.A2(net5),
.A3(in47),
.S0(net13),
.S1(net15),
.X(net21)
);

sky130_fd_sc_hd__and2_1 c84(
.A(net21),
.B(in58),
.X(net22)
);

sky130_fd_sc_hd__mux4_2 c85(
.A0(in28),
.A1(net18),
.A2(net21),
.A3(net5),
.S0(net12),
.S1(net6),
.X(net23)
);

sky130_fd_sc_hd__mux4_4 c86(
.A0(net17),
.A1(net21),
.A2(net23),
.A3(net22),
.S0(net20),
.S1(net2),
.X(net24)
);

sky130_fd_sc_hd__mux4_1 c87(
.A0(net18),
.A1(net24),
.A2(net23),
.A3(net22),
.S0(net5),
.S1(in28),
.X(net25)
);

sky130_fd_sc_hd__nor2b_4 c88(
.A(in20),
.B_N(in42),
.Y(net26)
);

sky130_fd_sc_hd__and2_4 c89(
.A(net15),
.B(net24),
.X(net27)
);

sky130_fd_sc_hd__nor2b_2 c90(
.A(in34),
.B_N(net15),
.Y(net28)
);

sky130_fd_sc_hd__a21boi_0 c91(
.A1(net22),
.A2(net16),
.B1_N(in51),
.Y(net29)
);

sky130_fd_sc_hd__mux4_4 c92(
.A0(in50),
.A1(net27),
.A2(net26),
.A3(in55),
.S0(net29),
.S1(net28),
.X(net30)
);

sky130_fd_sc_hd__nor2b_4 c93(
.A(in55),
.B_N(net7),
.Y(net31)
);

sky130_fd_sc_hd__and2_4 c94(
.A(in36),
.B(in3),
.X(net32)
);

sky130_fd_sc_hd__o21a_2 c95(
.A1(in51),
.A2(in34),
.B1(net26),
.X(net33)
);

sky130_fd_sc_hd__or2_1 c96(
.A(net29),
.B(net22),
.X(net34)
);

sky130_fd_sc_hd__nand2b_1 c97(
.A_N(net28),
.B(net33),
.Y(net35)
);

sky130_fd_sc_hd__and2b_4 c98(
.A_N(net35),
.B(net28),
.X(net36)
);

sky130_fd_sc_hd__a31oi_4 c99(
.A1(net34),
.A2(net30),
.A3(net15),
.B1(in59),
.Y(net37)
);

sky130_fd_sc_hd__nor2_2 c100(
.A(in30),
.B(net15),
.Y(net38)
);

sky130_fd_sc_hd__or2_4 c101(
.A(net36),
.B(in39),
.X(net39)
);

sky130_fd_sc_hd__and2b_4 c102(
.A_N(net27),
.B(in30),
.X(net40)
);

sky130_fd_sc_hd__a31o_1 c103(
.A1(net24),
.A2(net38),
.A3(net30),
.B1(net34),
.X(net41)
);

sky130_fd_sc_hd__mux4_4 c104(
.A0(net41),
.A1(net38),
.A2(in3),
.A3(net37),
.S0(net36),
.S1(net27),
.X(net42)
);

sky130_fd_sc_hd__a41oi_4 c105(
.A1(net39),
.A2(net38),
.A3(net41),
.A4(in49),
.B1(net22),
.Y(net43)
);

sky130_fd_sc_hd__mux2_4 c106(
.A0(net40),
.A1(net32),
.S(in50),
.X(net44)
);

sky130_fd_sc_hd__a31o_4 c107(
.A1(net44),
.A2(net27),
.A3(net38),
.B1(net29),
.X(net45)
);

sky130_fd_sc_hd__mux2_8 c108(
.A0(net36),
.A1(in44),
.S(net27),
.X(net46)
);

sky130_fd_sc_hd__a41oi_2 c109(
.A1(net46),
.A2(net26),
.A3(net37),
.A4(net35),
.B1(in59),
.Y(net47)
);

sky130_fd_sc_hd__nor2b_4 c110(
.A(net16),
.B_N(net42),
.Y(net48)
);

sky130_fd_sc_hd__nor2_1 c111(
.A(net17),
.B(net6),
.Y(net49)
);

sky130_fd_sc_hd__or2b_2 c112(
.A(net48),
.B_N(in13),
.X(net50)
);

sky130_fd_sc_hd__o21bai_1 c113(
.A1(in44),
.A2(in49),
.B1_N(in15),
.Y(net51)
);

sky130_fd_sc_hd__and2_2 c114(
.A(net47),
.B(net43),
.X(net52)
);

sky130_fd_sc_hd__nand2b_4 c115(
.A_N(net51),
.B(net47),
.Y(net53)
);

sky130_fd_sc_hd__nand2b_2 c116(
.A_N(net48),
.B(net32),
.Y(net54)
);

sky130_fd_sc_hd__or2_4 c117(
.A(net23),
.B(net52),
.X(net55)
);

sky130_fd_sc_hd__o21ai_1 c118(
.A1(net54),
.A2(net7),
.B1(net55),
.Y(net56)
);

sky130_fd_sc_hd__clkbuf_8 c119(
.A(net767),
.X(net57)
);

sky130_fd_sc_hd__a21o_2 c120(
.A1(net32),
.A2(net17),
.B1(net54),
.X(out57)
);

sky130_fd_sc_hd__mux4_2 c121(
.A0(in3),
.A1(net55),
.A2(net56),
.A3(net48),
.S0(net47),
.S1(net7),
.X(net58)
);

sky130_fd_sc_hd__buf_8 c122(
.A(net767),
.X(net59)
);

sky130_fd_sc_hd__nand2_4 c123(
.A(net57),
.B(net54),
.Y(net60)
);

sky130_fd_sc_hd__nand2b_2 c124(
.A_N(net53),
.B(net59),
.Y(net61)
);

sky130_fd_sc_hd__or2b_2 c125(
.A(net61),
.B_N(net29),
.X(net62)
);

sky130_fd_sc_hd__mux4_4 c126(
.A0(net60),
.A1(net61),
.A2(net50),
.A3(out57),
.S0(net54),
.S1(net790),
.X(net63)
);

sky130_fd_sc_hd__mux4_4 c127(
.A0(net11),
.A1(net62),
.A2(net60),
.A3(net47),
.S0(net789),
.S1(net791),
.X(net64)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c128(
.A(net767),
.X(net65)
);

sky130_fd_sc_hd__mux4_1 c129(
.A0(net65),
.A1(out57),
.A2(net42),
.A3(net54),
.S0(net59),
.S1(net792),
.X(net66)
);

sky130_fd_sc_hd__o21ai_2 c130(
.A1(net65),
.A2(net792),
.B1(net793),
.Y(net67)
);

sky130_fd_sc_hd__a21boi_1 c131(
.A1(net55),
.A2(net67),
.B1_N(net792),
.Y(net68)
);

sky130_fd_sc_hd__o21a_1 c132(
.A1(in18),
.A2(in11),
.B1(in14),
.X(net69)
);

sky130_fd_sc_hd__a31o_4 c133(
.A1(in17),
.A2(in1),
.A3(in19),
.B1(in7),
.X(net70)
);

sky130_fd_sc_hd__o21a_4 c134(
.A1(in4),
.A2(in2),
.B1(in8),
.X(net71)
);

sky130_fd_sc_hd__o21ai_2 c135(
.A1(in5),
.A2(net71),
.B1(in10),
.Y(net72)
);

sky130_fd_sc_hd__or2_1 c136(
.A(in6),
.B(in9),
.X(net73)
);

sky130_fd_sc_hd__and2b_1 c137(
.A_N(net71),
.B(in6),
.X(net74)
);

sky130_fd_sc_hd__nor2b_1 c138(
.A(in16),
.B_N(net74),
.Y(net75)
);

sky130_fd_sc_hd__a31o_4 c139(
.A1(net75),
.A2(in4),
.A3(in21),
.B1(in13),
.X(net76)
);

sky130_fd_sc_hd__nand2b_1 c140(
.A_N(in14),
.B(net75),
.Y(net77)
);

sky130_fd_sc_hd__o21ba_2 c141(
.A1(in21),
.A2(net72),
.B1_N(net75),
.X(net78)
);

sky130_fd_sc_hd__a31oi_1 c142(
.A1(net77),
.A2(in14),
.A3(in4),
.B1(net70),
.Y(net79)
);

sky130_fd_sc_hd__nand2b_1 c143(
.A_N(in5),
.B(in18),
.Y(net80)
);

sky130_fd_sc_hd__a31o_1 c144(
.A1(in2),
.A2(net76),
.A3(net73),
.B1(in13),
.X(net81)
);

sky130_fd_sc_hd__and2_0 c145(
.A(net75),
.B(net80),
.X(net82)
);

sky130_fd_sc_hd__nand2_1 c146(
.A(net82),
.B(net79),
.Y(net83)
);

sky130_fd_sc_hd__a31o_4 c147(
.A1(net81),
.A2(in1),
.A3(in6),
.B1(net75),
.X(net84)
);

sky130_fd_sc_hd__a41o_1 c148(
.A1(net83),
.A2(in0),
.A3(net74),
.A4(net76),
.B1(net84),
.X(net85)
);

sky130_fd_sc_hd__a41o_2 c149(
.A1(net80),
.A2(in21),
.A3(net77),
.A4(net75),
.B1(net83),
.X(net86)
);

sky130_fd_sc_hd__a31o_2 c150(
.A1(net70),
.A2(net78),
.A3(net82),
.B1(net69),
.X(net87)
);

sky130_fd_sc_hd__mux4_2 c151(
.A0(net84),
.A1(in16),
.A2(net82),
.A3(net77),
.S0(net85),
.S1(net83),
.X(net88)
);

sky130_fd_sc_hd__mux4_1 c152(
.A0(net86),
.A1(net78),
.A2(net84),
.A3(net87),
.S0(net83),
.S1(net70),
.X(net89)
);

sky130_fd_sc_hd__mux4_2 c153(
.A0(net88),
.A1(net89),
.A2(net81),
.A3(net73),
.S0(net86),
.S1(net78),
.X(net90)
);

sky130_fd_sc_hd__and2b_4 c154(
.A_N(in17),
.B(net88),
.X(net91)
);

sky130_fd_sc_hd__a21boi_1 c155(
.A1(in22),
.A2(in38),
.B1_N(in42),
.Y(net92)
);

sky130_fd_sc_hd__or2b_4 c156(
.A(net84),
.B_N(in35),
.X(net93)
);

sky130_fd_sc_hd__a41oi_1 c157(
.A1(in9),
.A2(in39),
.A3(net80),
.A4(net73),
.B1(net74),
.Y(net94)
);

sky130_fd_sc_hd__or2_2 c158(
.A(net78),
.B(in33),
.X(net95)
);

sky130_fd_sc_hd__o21ai_1 c159(
.A1(in1),
.A2(net94),
.B1(in22),
.Y(net96)
);

sky130_fd_sc_hd__and2b_2 c160(
.A_N(in23),
.B(in38),
.X(net97)
);

sky130_fd_sc_hd__or2b_2 c161(
.A(in27),
.B_N(net70),
.X(net98)
);

sky130_fd_sc_hd__nor2_4 c162(
.A(net95),
.B(net97),
.Y(net99)
);

sky130_fd_sc_hd__or2b_1 c163(
.A(net98),
.B_N(net99),
.X(net100)
);

sky130_fd_sc_hd__o21a_4 c164(
.A1(net88),
.A2(net92),
.B1(net97),
.X(net101)
);

sky130_fd_sc_hd__or2b_1 c165(
.A(net72),
.B_N(in42),
.X(net102)
);

sky130_fd_sc_hd__mux4_1 c166(
.A0(net97),
.A1(in15),
.A2(net96),
.A3(in29),
.S0(net102),
.S1(in39),
.X(net103)
);

sky130_fd_sc_hd__nor2_2 c167(
.A(in35),
.B(net93),
.Y(net104)
);

sky130_fd_sc_hd__a21oi_2 c168(
.A1(net102),
.A2(net89),
.B1(in23),
.Y(net105)
);

sky130_fd_sc_hd__a41o_4 c169(
.A1(net104),
.A2(net93),
.A3(in9),
.A4(in40),
.B1(net92),
.X(net106)
);

sky130_fd_sc_hd__a31o_2 c170(
.A1(in29),
.A2(net97),
.A3(net106),
.B1(in25),
.X(net107)
);

sky130_fd_sc_hd__a41o_1 c171(
.A1(in32),
.A2(net99),
.A3(net106),
.A4(net95),
.B1(net102),
.X(net108)
);

sky130_fd_sc_hd__a41o_2 c172(
.A1(net108),
.A2(net106),
.A3(net101),
.A4(net95),
.B1(net107),
.X(net109)
);

sky130_fd_sc_hd__mux4_1 c173(
.A0(net97),
.A1(net109),
.A2(net102),
.A3(in26),
.S0(net83),
.S1(net108),
.X(net110)
);

sky130_fd_sc_hd__mux4_1 c174(
.A0(net101),
.A1(net85),
.A2(net110),
.A3(in17),
.S0(in25),
.S1(net108),
.X(net111)
);

sky130_fd_sc_hd__a31o_4 c175(
.A1(net110),
.A2(in38),
.A3(net95),
.B1(net108),
.X(net112)
);

sky130_fd_sc_hd__nand2_4 c176(
.A(in26),
.B(in53),
.Y(net113)
);

sky130_fd_sc_hd__or2b_2 c177(
.A(net111),
.B_N(net3),
.X(net114)
);

sky130_fd_sc_hd__a31o_2 c178(
.A1(in60),
.A2(in19),
.A3(net114),
.B1(net110),
.X(net115)
);

sky130_fd_sc_hd__or2_4 c179(
.A(in12),
.B(net3),
.X(net116)
);

sky130_fd_sc_hd__or2b_1 c180(
.A(in25),
.B_N(net116),
.X(net117)
);

sky130_fd_sc_hd__a21oi_2 c181(
.A1(in52),
.A2(in46),
.B1(net99),
.Y(net118)
);

sky130_fd_sc_hd__and2b_2 c182(
.A_N(in48),
.B(net116),
.X(net119)
);

sky130_fd_sc_hd__a31o_2 c183(
.A1(net74),
.A2(net113),
.A3(in12),
.B1(net106),
.X(net120)
);

sky130_fd_sc_hd__nor2b_1 c184(
.A(net119),
.B_N(net106),
.Y(net121)
);

sky130_fd_sc_hd__a21bo_1 c185(
.A1(net117),
.A2(net116),
.B1_N(net121),
.X(net122)
);

sky130_fd_sc_hd__a21o_4 c186(
.A1(net118),
.A2(net73),
.B1(net122),
.X(net123)
);

sky130_fd_sc_hd__and2_4 c187(
.A(in57),
.B(net122),
.X(net124)
);

sky130_fd_sc_hd__mux4_2 c188(
.A0(in61),
.A1(net87),
.A2(net119),
.A3(net117),
.S0(net110),
.S1(in15),
.X(net125)
);

sky130_fd_sc_hd__a21boi_2 c189(
.A1(net123),
.A2(net122),
.B1_N(net125),
.Y(net126)
);

sky130_fd_sc_hd__a31o_4 c190(
.A1(net115),
.A2(net123),
.A3(net122),
.B1(net70),
.X(net127)
);

sky130_fd_sc_hd__a31o_1 c191(
.A1(net124),
.A2(in56),
.A3(net125),
.B1(net122),
.X(net128)
);

sky130_fd_sc_hd__clkbuf_2 c192(
.A(net721),
.X(net129)
);

sky130_fd_sc_hd__a31o_1 c193(
.A1(net73),
.A2(net128),
.A3(net122),
.B1(net722),
.X(net130)
);

sky130_fd_sc_hd__mux4_2 c194(
.A0(net114),
.A1(net118),
.A2(net129),
.A3(net122),
.S0(net124),
.S1(net123),
.X(out15)
);

sky130_fd_sc_hd__mux4_4 c195(
.A0(net129),
.A1(net126),
.A2(net122),
.A3(net99),
.S0(net114),
.S1(net721),
.X(net131)
);

sky130_fd_sc_hd__inv_16 c196(
.A(net721),
.Y(net132)
);

sky130_fd_sc_hd__mux4_1 c197(
.A0(net100),
.A1(in61),
.A2(net131),
.A3(net123),
.S0(net125),
.S1(net132),
.X(net133)
);

sky130_fd_sc_hd__and2_1 c198(
.A(net9),
.B(net110),
.X(net134)
);

sky130_fd_sc_hd__o21ai_1 c199(
.A1(net14),
.A2(net0),
.B1(net13),
.Y(net135)
);

sky130_fd_sc_hd__or2_2 c200(
.A(net135),
.B(net14),
.X(net136)
);

sky130_fd_sc_hd__mux2_2 c201(
.A0(net5),
.A1(net132),
.S(net1),
.X(net137)
);

sky130_fd_sc_hd__o21bai_1 c202(
.A1(net134),
.A2(net9),
.B1_N(net20),
.Y(net138)
);

sky130_fd_sc_hd__o21ai_2 c203(
.A1(in46),
.A2(net110),
.B1(net120),
.Y(net139)
);

sky130_fd_sc_hd__a41oi_1 c204(
.A1(net134),
.A2(net6),
.A3(net25),
.A4(net139),
.B1(net109),
.Y(net140)
);

sky130_fd_sc_hd__a21bo_2 c205(
.A1(net8),
.A2(net136),
.B1_N(net7),
.X(net141)
);

sky130_fd_sc_hd__mux2_2 c206(
.A0(net125),
.A1(net110),
.S(in42),
.X(net142)
);

sky130_fd_sc_hd__sdfrbp_1 c207(
.D(net132),
.RESET_B(net8),
.SCD(net142),
.SCE(net130),
.CLK(clk),
.Q(net144),
.Q_N(net143)
);

sky130_fd_sc_hd__a21oi_2 c208(
.A1(net136),
.A2(in8),
.B1(net7),
.Y(net145)
);

sky130_fd_sc_hd__nand2_4 c209(
.A(net142),
.B(in56),
.Y(net146)
);

sky130_fd_sc_hd__a31o_4 c210(
.A1(net141),
.A2(net83),
.A3(net145),
.B1(net114),
.X(net147)
);

sky130_fd_sc_hd__mux4_4 c211(
.A0(net13),
.A1(net135),
.A2(net132),
.A3(net143),
.S0(net147),
.S1(net141),
.X(net148)
);

sky130_fd_sc_hd__mux4_4 c212(
.A0(net135),
.A1(net140),
.A2(net83),
.A3(in46),
.S0(net147),
.S1(net737),
.X(net149)
);

sky130_fd_sc_hd__o21a_4 c213(
.A1(net4),
.A2(net142),
.B1(net736),
.X(net150)
);

sky130_fd_sc_hd__a41o_1 c214(
.A1(net144),
.A2(net99),
.A3(net150),
.A4(net147),
.B1(net736),
.X(net151)
);

sky130_fd_sc_hd__o21bai_2 c215(
.A1(net137),
.A2(in42),
.B1_N(in33),
.Y(net152)
);

sky130_fd_sc_hd__clkbuf_8 c216(
.A(net767),
.X(net153)
);

sky130_fd_sc_hd__a41o_2 c217(
.A1(net145),
.A2(net83),
.A3(net147),
.A4(net146),
.B1(net113),
.X(net154)
);

sky130_fd_sc_hd__mux4_2 c218(
.A0(net126),
.A1(net140),
.A2(net153),
.A3(net143),
.S0(in8),
.S1(net736),
.X(net155)
);

sky130_fd_sc_hd__a21oi_2 c219(
.A1(net152),
.A2(net99),
.B1(net751),
.Y(net156)
);

sky130_fd_sc_hd__nor2b_1 c220(
.A(net153),
.B_N(net137),
.Y(net157)
);

sky130_fd_sc_hd__or2b_4 c221(
.A(in38),
.B_N(net31),
.X(net158)
);

sky130_fd_sc_hd__a21oi_4 c222(
.A1(net157),
.A2(net137),
.B1(net794),
.Y(net159)
);

sky130_fd_sc_hd__and2b_1 c223(
.A_N(net109),
.B(net767),
.X(net160)
);

sky130_fd_sc_hd__and2b_4 c224(
.A_N(net28),
.B(net158),
.X(out55)
);

sky130_fd_sc_hd__nand2_4 c225(
.A(net159),
.B(net30),
.Y(net161)
);

sky130_fd_sc_hd__nand2_2 c226(
.A(net31),
.B(in59),
.Y(net162)
);

sky130_fd_sc_hd__a21boi_0 c227(
.A1(net120),
.A2(net137),
.B1_N(net29),
.Y(net163)
);

sky130_fd_sc_hd__mux4_2 c228(
.A0(net26),
.A1(net25),
.A2(in39),
.A3(out15),
.S0(net31),
.S1(net163),
.X(net164)
);

sky130_fd_sc_hd__nand2_4 c229(
.A(net138),
.B(net7),
.Y(net165)
);

sky130_fd_sc_hd__mux4_1 c230(
.A0(net37),
.A1(net43),
.A2(net159),
.A3(net7),
.S0(out55),
.S1(in39),
.X(net166)
);

sky130_fd_sc_hd__nand2_1 c231(
.A(net160),
.B(net162),
.Y(net167)
);

sky130_fd_sc_hd__mux4_2 c232(
.A0(net121),
.A1(net167),
.A2(net147),
.A3(net157),
.S0(net109),
.S1(net751),
.X(net168)
);

sky130_fd_sc_hd__a31o_4 c233(
.A1(net162),
.A2(in59),
.A3(net99),
.B1(out2),
.X(net169)
);

sky130_fd_sc_hd__mux4_4 c234(
.A0(net99),
.A1(in28),
.A2(net121),
.A3(net138),
.S0(net7),
.S1(net29),
.X(net170)
);

sky130_fd_sc_hd__clkinv_1 c235(
.A(net737),
.Y(net171)
);

sky130_fd_sc_hd__a31o_1 c236(
.A1(in59),
.A2(net169),
.A3(net767),
.B1(out2),
.X(net172)
);

sky130_fd_sc_hd__buf_8 c237(
.A(net737),
.X(net173)
);

sky130_fd_sc_hd__and2b_2 c238(
.A_N(net172),
.B(net138),
.X(net174)
);

sky130_fd_sc_hd__a31o_4 c239(
.A1(net30),
.A2(net172),
.A3(net105),
.B1(net169),
.X(net175)
);

sky130_fd_sc_hd__mux4_2 c240(
.A0(net174),
.A1(net137),
.A2(net170),
.A3(in53),
.S0(net25),
.S1(out2),
.X(net176)
);

sky130_fd_sc_hd__sdfbbn_1 c241(
.D(net175),
.RESET_B(net165),
.SCD(out15),
.SCE(net171),
.SET_B(net719),
.CLK_N(clk),
.Q(net178),
.Q_N(net177)
);

sky130_fd_sc_hd__a41oi_4 c242(
.A1(net50),
.A2(net49),
.A3(net719),
.A4(net722),
.B1(net790),
.Y(net179)
);

sky130_fd_sc_hd__a31oi_4 c243(
.A1(net52),
.A2(in56),
.A3(net751),
.B1(net790),
.Y(net180)
);

sky130_fd_sc_hd__a21o_1 c244(
.A1(net7),
.A2(net719),
.B1(net751),
.X(net181)
);

sky130_fd_sc_hd__mux2_2 c245(
.A0(net166),
.A1(net50),
.S(net109),
.X(net182)
);

sky130_fd_sc_hd__inv_16 c246(
.A(net697),
.Y(net183)
);

sky130_fd_sc_hd__o21bai_4 c247(
.A1(net52),
.A2(net181),
.B1_N(net789),
.Y(net184)
);

sky130_fd_sc_hd__clkbuf_4 c248(
.A(net697),
.X(out28)
);

sky130_fd_sc_hd__a31o_1 c249(
.A1(net180),
.A2(net6),
.A3(net177),
.B1(in42),
.X(net185)
);

sky130_fd_sc_hd__clkinv_4 c250(
.A(net767),
.Y(out27)
);

sky130_fd_sc_hd__o21bai_2 c251(
.A1(net49),
.A2(in42),
.B1_N(net184),
.Y(net186)
);

sky130_fd_sc_hd__o21ai_0 c252(
.A1(net183),
.A2(net185),
.B1(net68),
.Y(net187)
);

sky130_fd_sc_hd__inv_16 c253(
.A(net767),
.Y(out60)
);

sky130_fd_sc_hd__a31o_4 c254(
.A1(net181),
.A2(out60),
.A3(net184),
.B1(out49),
.X(net188)
);

sky130_fd_sc_hd__mux4_2 c255(
.A0(net43),
.A1(out57),
.A2(out60),
.A3(net178),
.S0(net49),
.S1(out55),
.X(net189)
);

sky130_fd_sc_hd__buf_16 c256(
.A(net719),
.X(net190)
);

sky130_fd_sc_hd__sdfbbn_2 c257(
.D(net50),
.RESET_B(net188),
.SCD(net33),
.SCE(net793),
.SET_B(net795),
.CLK_N(clk),
.Q(net192),
.Q_N(net191)
);

sky130_fd_sc_hd__o21ba_1 c258(
.A1(net184),
.A2(net109),
.B1_N(net795),
.X(net193)
);

sky130_fd_sc_hd__a21boi_2 c259(
.A1(net192),
.A2(out60),
.B1_N(net722),
.Y(net194)
);

sky130_fd_sc_hd__mux4_2 c260(
.A0(net186),
.A1(net194),
.A2(net50),
.A3(net188),
.S0(net49),
.S1(out55),
.X(net195)
);

sky130_fd_sc_hd__mux4_1 c261(
.A0(in15),
.A1(net194),
.A2(net192),
.A3(net43),
.S0(net188),
.S1(net751),
.X(net196)
);

sky130_fd_sc_hd__sdfbbp_1 c262(
.D(net171),
.RESET_B(net193),
.SCD(net191),
.SCE(net751),
.SET_B(net796),
.CLK(clk),
.Q(net198),
.Q_N(net197)
);

sky130_fd_sc_hd__mux4_2 c263(
.A0(net190),
.A1(net191),
.A2(net197),
.A3(net751),
.S0(out2),
.S1(net796),
.X(net199)
);

sky130_fd_sc_hd__a21o_2 c264(
.A1(net72),
.A2(net73),
.B1(net87),
.X(net200)
);

sky130_fd_sc_hd__nor2_1 c265(
.A(net82),
.B(net90),
.Y(net201)
);

sky130_fd_sc_hd__and2b_4 c266(
.A_N(net76),
.B(net90),
.X(net202)
);

sky130_fd_sc_hd__and2b_4 c267(
.A_N(net202),
.B(net87),
.X(net203)
);

sky130_fd_sc_hd__nand2_2 c268(
.A(net202),
.B(net85),
.Y(net204)
);

sky130_fd_sc_hd__a21bo_1 c269(
.A1(net203),
.A2(net87),
.B1_N(net77),
.X(net205)
);

sky130_fd_sc_hd__or2b_4 c270(
.A(net200),
.B_N(net202),
.X(net206)
);

sky130_fd_sc_hd__nand2_1 c271(
.A(net87),
.B(net203),
.Y(net207)
);

sky130_fd_sc_hd__nand2_4 c272(
.A(net205),
.B(net204),
.Y(net208)
);

sky130_fd_sc_hd__xor2_2 c273(
.A(net202),
.B(net90),
.X(net209)
);

sky130_fd_sc_hd__xnor2_4 c274(
.A(net204),
.B(net208),
.Y(net210)
);

sky130_fd_sc_hd__a21bo_1 c275(
.A1(net207),
.A2(in10),
.B1_N(net202),
.X(net211)
);

sky130_fd_sc_hd__xor2_1 c276(
.A(net208),
.B(in10),
.X(net212)
);

sky130_fd_sc_hd__o21bai_4 c277(
.A1(net212),
.A2(net202),
.B1_N(in4),
.Y(net213)
);

sky130_fd_sc_hd__clkinv_4 c278(
.A(net703),
.Y(net214)
);

sky130_fd_sc_hd__mux4_2 c279(
.A0(net213),
.A1(net71),
.A2(net214),
.A3(in8),
.S0(net205),
.S1(net203),
.X(net215)
);

sky130_fd_sc_hd__mux4_1 c280(
.A0(net85),
.A1(net213),
.A2(net204),
.A3(in14),
.S0(net205),
.S1(net69),
.X(net216)
);

sky130_fd_sc_hd__a21oi_4 c281(
.A1(in11),
.A2(net703),
.B1(net798),
.Y(net217)
);

sky130_fd_sc_hd__xor2_2 c282(
.A(net209),
.B(net798),
.X(net218)
);

sky130_fd_sc_hd__a31o_4 c283(
.A1(net210),
.A2(net212),
.A3(net217),
.B1(net703),
.X(net219)
);

sky130_fd_sc_hd__inv_2 c284(
.A(net703),
.Y(net220)
);

sky130_fd_sc_hd__mux4_1 c285(
.A0(net219),
.A1(net220),
.A2(net217),
.A3(net212),
.S0(net213),
.S1(net703),
.X(net221)
);

sky130_fd_sc_hd__xnor2_4 c286(
.A(net210),
.B(net72),
.Y(out33)
);

sky130_fd_sc_hd__o21bai_2 c287(
.A1(net91),
.A2(net94),
.B1_N(in39),
.Y(net222)
);

sky130_fd_sc_hd__a31oi_1 c288(
.A1(net208),
.A2(net200),
.A3(net83),
.B1(net81),
.Y(net223)
);

sky130_fd_sc_hd__a41oi_4 c289(
.A1(net222),
.A2(net94),
.A3(net210),
.A4(net206),
.B1(net203),
.Y(net224)
);

sky130_fd_sc_hd__inv_8 c290(
.A(net781),
.Y(net225)
);

sky130_fd_sc_hd__xor2_2 c291(
.A(net109),
.B(net206),
.X(net226)
);

sky130_fd_sc_hd__xor2_1 c292(
.A(net94),
.B(in10),
.X(net227)
);

sky130_fd_sc_hd__o21ba_2 c293(
.A1(in37),
.A2(net223),
.B1_N(net108),
.X(net228)
);

sky130_fd_sc_hd__xnor2_1 c294(
.A(in40),
.B(net205),
.Y(out8)
);

sky130_fd_sc_hd__buf_12 c295(
.A(net781),
.X(net229)
);

sky130_fd_sc_hd__mux4_4 c296(
.A0(net229),
.A1(net227),
.A2(in37),
.A3(net87),
.S0(net222),
.S1(net224),
.X(net230)
);

sky130_fd_sc_hd__sdfbbn_1 c297(
.D(net89),
.RESET_B(net228),
.SCD(net94),
.SCE(in8),
.SET_B(net797),
.CLK_N(clk),
.Q(net232),
.Q_N(net231)
);

sky130_fd_sc_hd__xor2_4 c298(
.A(net103),
.B(out8),
.X(net233)
);

sky130_fd_sc_hd__o21ai_0 c299(
.A1(in31),
.A2(net223),
.B1(out8),
.Y(net234)
);

sky130_fd_sc_hd__xor2_2 c300(
.A(net206),
.B(net227),
.X(net235)
);

sky130_fd_sc_hd__mux2_1 c301(
.A0(net96),
.A1(net214),
.S(out8),
.X(net236)
);

sky130_fd_sc_hd__mux4_2 c302(
.A0(net232),
.A1(net234),
.A2(net224),
.A3(net228),
.S0(net93),
.S1(out33),
.X(net237)
);

sky130_fd_sc_hd__a41oi_4 c303(
.A1(net112),
.A2(net210),
.A3(net234),
.A4(net94),
.B1(net235),
.Y(net238)
);

sky130_fd_sc_hd__a21o_4 c304(
.A1(net235),
.A2(net203),
.B1(net781),
.X(net239)
);

sky130_fd_sc_hd__sdfbbn_2 c305(
.D(net234),
.RESET_B(net239),
.SCD(net229),
.SCE(out8),
.SET_B(net781),
.CLK_N(clk),
.Q(net241),
.Q_N(net240)
);

sky130_fd_sc_hd__a41oi_2 c306(
.A1(net241),
.A2(out8),
.A3(net235),
.A4(net223),
.B1(net742),
.Y(out18)
);

sky130_fd_sc_hd__mux4_2 c307(
.A0(net233),
.A1(net232),
.A2(net239),
.A3(net234),
.S0(net89),
.S1(net240),
.X(net242)
);

sky130_fd_sc_hd__xnor2_1 c308(
.A(net200),
.B(in54),
.Y(net243)
);

sky130_fd_sc_hd__clkbuf_8 c309(
.A(net764),
.X(net244)
);

sky130_fd_sc_hd__dlygate4sd3_1 c310(
.A(net783),
.X(net245)
);

sky130_fd_sc_hd__o21bai_1 c311(
.A1(net245),
.A2(net107),
.B1_N(net226),
.Y(net246)
);

sky130_fd_sc_hd__inv_16 c312(
.A(net764),
.Y(net247)
);

sky130_fd_sc_hd__o21bai_2 c313(
.A1(net202),
.A2(net109),
.B1_N(net247),
.Y(net248)
);

sky130_fd_sc_hd__inv_4 c314(
.A(net742),
.Y(net249)
);

sky130_fd_sc_hd__xnor2_2 c315(
.A(net244),
.B(net122),
.Y(net250)
);

sky130_fd_sc_hd__xor2_1 c316(
.A(net249),
.B(net247),
.X(net251)
);

sky130_fd_sc_hd__mux4_2 c317(
.A0(net246),
.A1(net130),
.A2(net251),
.A3(net227),
.S0(net741),
.S1(net781),
.X(net252)
);

sky130_fd_sc_hd__mux4_2 c318(
.A0(in54),
.A1(net248),
.A2(net107),
.A3(net246),
.S0(net1),
.S1(net774),
.X(net253)
);

sky130_fd_sc_hd__mux2_8 c319(
.A0(net123),
.A1(net227),
.S(net253),
.X(net254)
);

sky130_fd_sc_hd__a41oi_4 c320(
.A1(net250),
.A2(net245),
.A3(net254),
.A4(net202),
.B1(net108),
.Y(net255)
);

sky130_fd_sc_hd__mux4_4 c321(
.A0(net122),
.A1(in53),
.A2(net105),
.A3(net253),
.S0(net106),
.S1(net80),
.X(net256)
);

sky130_fd_sc_hd__buf_8 c322(
.A(net783),
.X(net257)
);

sky130_fd_sc_hd__dlygate4sd1_1 c323(
.A(net745),
.X(net258)
);

sky130_fd_sc_hd__xnor2_4 c324(
.A(net251),
.B(net257),
.Y(net259)
);

sky130_fd_sc_hd__mux4_1 c325(
.A0(net258),
.A1(net250),
.A2(net256),
.A3(net128),
.S0(net123),
.S1(net259),
.X(net260)
);

sky130_fd_sc_hd__mux4_2 c326(
.A0(net254),
.A1(net123),
.A2(net259),
.A3(net246),
.S0(net741),
.S1(net783),
.X(net261)
);

sky130_fd_sc_hd__mux4_1 c327(
.A0(net249),
.A1(net258),
.A2(net254),
.A3(in42),
.S0(net783),
.S1(net800),
.X(net262)
);

sky130_fd_sc_hd__a41oi_2 c328(
.A1(net243),
.A2(net259),
.A3(net244),
.A4(net774),
.B1(net783),
.Y(net263)
);

sky130_fd_sc_hd__sdfbbp_1 c329(
.D(net253),
.RESET_B(net228),
.SCD(net755),
.SCE(net781),
.SET_B(net783),
.CLK(clk),
.Q(out38),
.Q_N(net264)
);

sky130_fd_sc_hd__xor2_2 c330(
.A(net251),
.B(net232),
.X(net265)
);

sky130_fd_sc_hd__a21boi_2 c331(
.A1(net265),
.A2(net755),
.B1_N(net799),
.Y(net266)
);

sky130_fd_sc_hd__a21o_1 c332(
.A1(net128),
.A2(net220),
.B1(net799),
.X(net267)
);

sky130_fd_sc_hd__sdfbbn_1 c333(
.D(net266),
.RESET_B(net140),
.SCD(net267),
.SCE(net114),
.SET_B(net781),
.CLK_N(clk),
.Q(out26),
.Q_N(net268)
);

sky130_fd_sc_hd__sdfrbp_2 c334(
.D(net150),
.RESET_B(net2),
.SCD(net155),
.SCE(net114),
.CLK(clk),
.Q(net270),
.Q_N(net269)
);

sky130_fd_sc_hd__xor2_1 c335(
.A(net156),
.B(in39),
.X(net271)
);

sky130_fd_sc_hd__xor2_4 c336(
.A(net83),
.B(net269),
.X(net272)
);

sky130_fd_sc_hd__mux4_4 c337(
.A0(net114),
.A1(net25),
.A2(net128),
.A3(net156),
.S0(net272),
.S1(net271),
.X(net273)
);

sky130_fd_sc_hd__buf_8 c338(
.A(net765),
.X(net274)
);

sky130_fd_sc_hd__inv_12 c339(
.A(net764),
.Y(net275)
);

sky130_fd_sc_hd__a41oi_2 c340(
.A1(net270),
.A2(net225),
.A3(net19),
.A4(net794),
.B1(net799),
.Y(net276)
);

sky130_fd_sc_hd__xnor2_4 c341(
.A(net220),
.B(net275),
.Y(net277)
);

sky130_fd_sc_hd__o21ai_4 c342(
.A1(net20),
.A2(net225),
.B1(net277),
.Y(net278)
);

sky130_fd_sc_hd__xor2_2 c343(
.A(net277),
.B(net755),
.X(out43)
);

sky130_fd_sc_hd__a41o_4 c344(
.A1(net225),
.A2(net270),
.A3(net276),
.A4(net278),
.B1(net774),
.X(net279)
);

sky130_fd_sc_hd__mux4_4 c345(
.A0(net248),
.A1(net83),
.A2(net265),
.A3(net267),
.S0(net278),
.S1(net266),
.X(net280)
);

sky130_fd_sc_hd__xnor2_1 c346(
.A(net277),
.B(net144),
.Y(net281)
);

sky130_fd_sc_hd__mux4_2 c347(
.A0(net257),
.A1(net281),
.A2(net150),
.A3(out8),
.S0(net278),
.S1(net225),
.X(net282)
);

sky130_fd_sc_hd__mux4_1 c348(
.A0(net279),
.A1(net20),
.A2(net272),
.A3(net267),
.S0(net278),
.S1(out44),
.X(net283)
);

sky130_fd_sc_hd__mux4_2 c349(
.A0(net6),
.A1(net277),
.A2(net113),
.A3(net278),
.S0(net273),
.S1(net729),
.X(net284)
);

sky130_fd_sc_hd__mux4_1 c350(
.A0(net277),
.A1(net279),
.A2(net267),
.A3(out43),
.S0(net278),
.S1(out44),
.X(net285)
);

sky130_fd_sc_hd__mux4_4 c351(
.A0(net144),
.A1(out26),
.A2(net231),
.A3(net729),
.S0(net757),
.S1(out44),
.X(net286)
);

sky130_fd_sc_hd__a31o_4 c352(
.A1(net173),
.A2(in7),
.A3(net271),
.B1(net33),
.X(net287)
);

sky130_fd_sc_hd__a31o_2 c353(
.A1(net147),
.A2(net140),
.A3(net281),
.B1(net774),
.X(net288)
);

sky130_fd_sc_hd__xor2_2 c354(
.A(net276),
.B(net278),
.X(net289)
);

sky130_fd_sc_hd__a31o_1 c355(
.A1(net281),
.A2(net163),
.A3(net278),
.B1(net800),
.X(net290)
);

sky130_fd_sc_hd__a31o_4 c356(
.A1(net271),
.A2(net161),
.A3(net231),
.B1(net800),
.X(out45)
);

sky130_fd_sc_hd__o21a_2 c357(
.A1(in53),
.A2(out45),
.B1(net278),
.X(net291)
);

sky130_fd_sc_hd__xnor2_2 c358(
.A(net278),
.B(out43),
.Y(net292)
);

sky130_fd_sc_hd__sdfbbn_2 c359(
.D(net147),
.RESET_B(net292),
.SCD(net140),
.SCE(net794),
.SET_B(out2),
.CLK_N(clk),
.Q(net294),
.Q_N(net293)
);

sky130_fd_sc_hd__mux4_4 c360(
.A0(net289),
.A1(net292),
.A2(net6),
.A3(net293),
.S0(net109),
.S1(net291),
.X(net295)
);

sky130_fd_sc_hd__a31o_2 c361(
.A1(net286),
.A2(net12),
.A3(net276),
.B1(in7),
.X(net296)
);

sky130_fd_sc_hd__mux4_1 c362(
.A0(net232),
.A1(in56),
.A2(net42),
.A3(net292),
.S0(out55),
.S1(net293),
.X(net297)
);

sky130_fd_sc_hd__a31o_1 c363(
.A1(net296),
.A2(net147),
.A3(net38),
.B1(net757),
.X(net298)
);

sky130_fd_sc_hd__sdfbbp_1 c364(
.D(net140),
.RESET_B(out33),
.SCD(net292),
.SCE(net6),
.SET_B(net794),
.CLK(clk),
.Q(out37),
.Q_N(net299)
);

sky130_fd_sc_hd__a41oi_1 c365(
.A1(net294),
.A2(net139),
.A3(net292),
.A4(net299),
.B1(net800),
.Y(net300)
);

sky130_fd_sc_hd__a41o_4 c366(
.A1(net297),
.A2(out43),
.A3(net173),
.A4(net299),
.B1(net757),
.X(net301)
);

sky130_fd_sc_hd__mux4_1 c367(
.A0(net301),
.A1(in7),
.A2(net231),
.A3(net33),
.S0(net294),
.S1(net299),
.X(net302)
);

sky130_fd_sc_hd__clkbuf_8 c368(
.A(net719),
.X(net303)
);

sky130_fd_sc_hd__a41oi_4 c369(
.A1(net295),
.A2(net296),
.A3(net302),
.A4(net303),
.B1(net299),
.Y(net304)
);

sky130_fd_sc_hd__mux4_2 c370(
.A0(net292),
.A1(net301),
.A2(net289),
.A3(in49),
.S0(out55),
.S1(net147),
.X(net305)
);

sky130_fd_sc_hd__mux4_4 c371(
.A0(net286),
.A1(out45),
.A2(in49),
.A3(net302),
.S0(net299),
.S1(net765),
.X(net306)
);

sky130_fd_sc_hd__a41oi_2 c372(
.A1(net271),
.A2(net292),
.A3(net299),
.A4(out42),
.B1(net765),
.Y(net307)
);

sky130_fd_sc_hd__mux4_4 c373(
.A0(net307),
.A1(net296),
.A2(in56),
.A3(net299),
.S0(net765),
.S1(net773),
.X(net308)
);

sky130_fd_sc_hd__clkbuf_4 c374(
.A(out20),
.X(net309)
);

sky130_fd_sc_hd__mux4_2 c375(
.A0(net309),
.A1(out57),
.A2(out27),
.A3(net68),
.S0(net299),
.S1(net795),
.X(net310)
);

sky130_fd_sc_hd__o21bai_4 c376(
.A1(net192),
.A2(net109),
.B1_N(net309),
.Y(out52)
);

sky130_fd_sc_hd__a21oi_1 c377(
.A1(out42),
.A2(net793),
.B1(out34),
.Y(net311)
);

sky130_fd_sc_hd__buf_4 c378(
.A(out20),
.X(net312)
);

sky130_fd_sc_hd__a41o_2 c379(
.A1(net68),
.A2(net309),
.A3(net199),
.A4(net773),
.B1(out2),
.X(net313)
);

sky130_fd_sc_hd__o21ba_1 c380(
.A1(net139),
.A2(in42),
.B1_N(net773),
.X(net314)
);

sky130_fd_sc_hd__a41oi_2 c381(
.A1(in42),
.A2(net300),
.A3(net33),
.A4(out42),
.B1(out53),
.Y(net315)
);

sky130_fd_sc_hd__a41o_1 c382(
.A1(net300),
.A2(net198),
.A3(out60),
.A4(out52),
.B1(net796),
.X(net316)
);

sky130_fd_sc_hd__mux4_1 c383(
.A0(net178),
.A1(net316),
.A2(net314),
.A3(net197),
.S0(out34),
.S1(net795),
.X(net317)
);

sky130_fd_sc_hd__mux4_4 c384(
.A0(in56),
.A1(net198),
.A2(net139),
.A3(net316),
.S0(net33),
.S1(net773),
.X(net318)
);

sky130_fd_sc_hd__mux4_4 c385(
.A0(net42),
.A1(net314),
.A2(net199),
.A3(net177),
.S0(net264),
.S1(net795),
.X(out14)
);

sky130_fd_sc_hd__clkinv_16 c386(
.A(net745),
.Y(out50)
);

sky130_fd_sc_hd__a41oi_1 c387(
.A1(net302),
.A2(out52),
.A3(net139),
.A4(net316),
.B1(in56),
.Y(net319)
);

sky130_fd_sc_hd__buf_4 c388(
.A(net788),
.X(out46)
);

sky130_fd_sc_hd__a41o_2 c389(
.A1(net33),
.A2(net314),
.A3(out52),
.A4(out46),
.B1(out55),
.X(net320)
);

sky130_fd_sc_hd__mux4_1 c390(
.A0(net312),
.A1(net198),
.A2(out37),
.A3(net290),
.S0(in56),
.S1(net268),
.X(out58)
);

sky130_fd_sc_hd__a31oi_2 c391(
.A1(net316),
.A2(out33),
.A3(net290),
.B1(net763),
.Y(net321)
);

sky130_fd_sc_hd__a41oi_1 c392(
.A1(net290),
.A2(out46),
.A3(net264),
.A4(net793),
.B1(out34),
.Y(out56)
);

sky130_fd_sc_hd__mux4_4 c393(
.A0(net314),
.A1(out28),
.A2(out56),
.A3(net139),
.S0(out46),
.S1(net793),
.X(net322)
);

sky130_fd_sc_hd__mux4_2 c394(
.A0(net322),
.A1(net316),
.A2(out56),
.A3(out46),
.S0(out37),
.S1(out22),
.X(net323)
);

sky130_fd_sc_hd__a41oi_1 c395(
.A1(net320),
.A2(net316),
.A3(net139),
.A4(net763),
.B1(out20),
.Y(net324)
);

sky130_fd_sc_hd__xnor2_4 c396(
.A(net212),
.B(net71),
.Y(net325)
);

sky130_fd_sc_hd__inv_6 c397(
.A(net718),
.Y(net326)
);

sky130_fd_sc_hd__a21bo_2 c398(
.A1(net71),
.A2(in8),
.B1_N(net797),
.X(net327)
);

sky130_fd_sc_hd__o21ai_0 c399(
.A1(net79),
.A2(net211),
.B1(in14),
.Y(net328)
);

sky130_fd_sc_hd__xnor2_1 c400(
.A(net76),
.B(net71),
.Y(net329)
);

sky130_fd_sc_hd__xor2_4 c401(
.A(net327),
.B(net211),
.X(net330)
);

sky130_fd_sc_hd__a31oi_2 c402(
.A1(net73),
.A2(net330),
.A3(net218),
.B1(net209),
.Y(net331)
);

sky130_fd_sc_hd__o21a_4 c403(
.A1(net326),
.A2(net212),
.B1(net209),
.X(net332)
);

sky130_fd_sc_hd__xnor2_2 c404(
.A(in11),
.B(in0),
.Y(net333)
);

sky130_fd_sc_hd__xnor2_2 c405(
.A(net328),
.B(net69),
.Y(net334)
);

sky130_fd_sc_hd__buf_12 c406(
.A(net694),
.X(net335)
);

sky130_fd_sc_hd__buf_8 c407(
.A(net694),
.X(net336)
);

sky130_fd_sc_hd__mux4_2 c408(
.A0(net325),
.A1(net336),
.A2(net334),
.A3(net326),
.S0(net329),
.S1(net330),
.X(net337)
);

sky130_fd_sc_hd__mux4_4 c409(
.A0(net336),
.A1(net327),
.A2(net218),
.A3(net334),
.S0(net326),
.S1(net330),
.X(net338)
);

sky130_fd_sc_hd__o21ai_4 c410(
.A1(net333),
.A2(net326),
.B1(net335),
.Y(net339)
);

sky130_fd_sc_hd__o21ai_4 c411(
.A1(net339),
.A2(net336),
.B1(net802),
.Y(net340)
);

sky130_fd_sc_hd__a31oi_4 c412(
.A1(net326),
.A2(net335),
.A3(net339),
.B1(net695),
.Y(net341)
);

sky130_fd_sc_hd__o21a_2 c413(
.A1(net335),
.A2(net339),
.B1(net802),
.X(net342)
);

sky130_fd_sc_hd__sdfbbn_1 c414(
.D(net341),
.RESET_B(net325),
.SCD(net339),
.SCE(net69),
.SET_B(net801),
.CLK_N(clk),
.Q(net344),
.Q_N(net343)
);

sky130_fd_sc_hd__mux2_1 c415(
.A0(net69),
.A1(net339),
.S(net341),
.X(net345)
);

sky130_fd_sc_hd__mux4_1 c416(
.A0(net345),
.A1(net341),
.A2(net339),
.A3(net336),
.S0(net344),
.S1(net330),
.X(net346)
);

sky130_fd_sc_hd__inv_8 c417(
.A(net718),
.Y(net347)
);

sky130_fd_sc_hd__clkinv_8 c418(
.A(net740),
.Y(net348)
);

sky130_fd_sc_hd__inv_6 c419(
.A(net740),
.Y(net349)
);

sky130_fd_sc_hd__sdfbbn_2 c420(
.D(net349),
.RESET_B(net330),
.SCD(net205),
.SCE(net331),
.SET_B(net348),
.CLK_N(clk),
.Q(net351),
.Q_N(net350)
);

sky130_fd_sc_hd__o21ba_2 c421(
.A1(net205),
.A2(net241),
.B1_N(net344),
.X(net352)
);

sky130_fd_sc_hd__o21ai_1 c422(
.A1(in0),
.A2(net227),
.B1(net798),
.Y(net353)
);

sky130_fd_sc_hd__a41oi_4 c423(
.A1(net92),
.A2(net342),
.A3(net240),
.A4(out18),
.B1(net801),
.Y(net354)
);

sky130_fd_sc_hd__mux2_2 c424(
.A0(net203),
.A1(net205),
.S(net755),
.X(net355)
);

sky130_fd_sc_hd__mux2_4 c425(
.A0(net355),
.A1(net348),
.S(net798),
.X(net356)
);

sky130_fd_sc_hd__a31o_2 c426(
.A1(net241),
.A2(net353),
.A3(net107),
.B1(net350),
.X(net357)
);

sky130_fd_sc_hd__o21bai_4 c427(
.A1(net357),
.A2(net348),
.B1_N(net343),
.Y(net358)
);

sky130_fd_sc_hd__mux2_8 c428(
.A0(net353),
.A1(net356),
.S(net358),
.X(net359)
);

sky130_fd_sc_hd__a21bo_4 c429(
.A1(net352),
.A2(net240),
.B1_N(net358),
.X(net360)
);

sky130_fd_sc_hd__inv_2 c430(
.A(net739),
.Y(net361)
);

sky130_fd_sc_hd__a21oi_4 c431(
.A1(net360),
.A2(net358),
.B1(net361),
.Y(net362)
);

sky130_fd_sc_hd__sdfrtn_1 c432(
.D(net361),
.RESET_B(net362),
.SCD(net348),
.SCE(net350),
.CLK_N(clk),
.Q(net363)
);

sky130_fd_sc_hd__buf_12 c433(
.A(net747),
.X(net364)
);

sky130_fd_sc_hd__a21boi_0 c434(
.A1(net355),
.A2(net357),
.B1_N(net364),
.Y(net365)
);

sky130_fd_sc_hd__clkbuf_16 c435(
.A(net779),
.X(net366)
);

sky130_fd_sc_hd__mux4_4 c436(
.A0(in41),
.A1(net355),
.A2(net364),
.A3(net366),
.S0(in39),
.S1(net92),
.X(net367)
);

sky130_fd_sc_hd__mux4_4 c437(
.A0(net364),
.A1(net367),
.A2(net366),
.A3(net363),
.S0(net355),
.S1(net344),
.X(net368)
);

sky130_fd_sc_hd__inv_2 c438(
.A(net747),
.Y(net369)
);

sky130_fd_sc_hd__mux4_4 c439(
.A0(net362),
.A1(net369),
.A2(net368),
.A3(net367),
.S0(net342),
.S1(net802),
.X(net370)
);

sky130_fd_sc_hd__clkinv_8 c440(
.A(net743),
.Y(out54)
);

sky130_fd_sc_hd__xnor2_2 c441(
.A(net107),
.B(in33),
.Y(net371)
);

sky130_fd_sc_hd__xnor2_1 c442(
.A(net239),
.B(net794),
.Y(net372)
);

sky130_fd_sc_hd__xnor2_1 c443(
.A(net203),
.B(net371),
.Y(out7)
);

sky130_fd_sc_hd__a41oi_1 c444(
.A1(out54),
.A2(net366),
.A3(net203),
.A4(net794),
.B1(net799),
.Y(net373)
);

sky130_fd_sc_hd__buf_2 c445(
.A(net743),
.X(net374)
);

sky130_fd_sc_hd__xnor2_4 c446(
.A(net372),
.B(net366),
.Y(net375)
);

sky130_fd_sc_hd__mux4_2 c447(
.A0(net365),
.A1(net239),
.A2(net253),
.A3(net375),
.S0(net254),
.S1(net794),
.X(net376)
);

sky130_fd_sc_hd__o21ai_4 c448(
.A1(net80),
.A2(in33),
.B1(net246),
.Y(net377)
);

sky130_fd_sc_hd__a41o_2 c449(
.A1(net371),
.A2(net377),
.A3(net348),
.A4(net342),
.B1(net794),
.X(net378)
);

sky130_fd_sc_hd__xor2_4 c450(
.A(net356),
.B(net246),
.X(net379)
);

sky130_fd_sc_hd__a41oi_4 c451(
.A1(net106),
.A2(net378),
.A3(net379),
.A4(out7),
.B1(net130),
.Y(net380)
);

sky130_fd_sc_hd__mux4_1 c452(
.A0(net378),
.A1(out54),
.A2(net379),
.A3(net203),
.S0(in33),
.S1(net263),
.X(net381)
);

sky130_fd_sc_hd__mux4_2 c453(
.A0(net227),
.A1(net70),
.A2(net363),
.A3(net379),
.S0(in7),
.S1(net803),
.X(net382)
);

sky130_fd_sc_hd__mux4_2 c454(
.A0(net375),
.A1(out54),
.A2(net373),
.A3(net348),
.S0(net803),
.S1(net804),
.X(net383)
);

sky130_fd_sc_hd__mux4_1 c455(
.A0(net263),
.A1(net246),
.A2(net113),
.A3(net253),
.S0(net804),
.S1(net805),
.X(net384)
);

sky130_fd_sc_hd__buf_1 c456(
.A(net745),
.X(net385)
);

sky130_fd_sc_hd__mux4_2 c457(
.A0(net253),
.A1(net106),
.A2(out7),
.A3(net365),
.S0(net348),
.S1(net342),
.X(net386)
);

sky130_fd_sc_hd__mux4_1 c458(
.A0(net377),
.A1(net342),
.A2(net366),
.A3(net384),
.S0(net803),
.S1(net805),
.X(net387)
);

sky130_fd_sc_hd__mux4_1 c459(
.A0(net1),
.A1(net113),
.A2(net253),
.A3(net386),
.S0(net733),
.X(net388)
);

sky130_fd_sc_hd__mux4_1 c460(
.A0(net386),
.A1(net379),
.A2(net254),
.A3(net108),
.S0(net733),
.S1(net804),
.X(net389)
);

sky130_fd_sc_hd__mux4_4 c461(
.A0(net253),
.A1(out54),
.A2(net748),
.A3(net803),
.S0(net805),
.S1(net806),
.X(net390)
);

sky130_fd_sc_hd__sdfbbp_1 c462(
.D(net342),
.RESET_B(out41),
.SCD(in39),
.SCE(net273),
.SET_B(net804),
.CLK(clk),
.Q(net392),
.Q_N(net391)
);

sky130_fd_sc_hd__a41oi_2 c463(
.A1(net406),
.A2(net363),
.A3(net348),
.A4(in19),
.B1(net269),
.Y(net393)
);

sky130_fd_sc_hd__mux4_2 c464(
.A0(net407),
.A1(net408),
.A2(net108),
.A3(out43),
.S0(net781),
.S1(net804),
.X(net394)
);

sky130_fd_sc_hd__a21boi_4 c465(
.A1(in8),
.A2(net259),
.B1_N(net407),
.Y(net395)
);

sky130_fd_sc_hd__mux2_2 c466(
.A0(net275),
.A1(net395),
.S(net410),
.X(net396)
);

sky130_fd_sc_hd__a41oi_2 c467(
.A1(net363),
.A2(net407),
.A3(out54),
.A4(net1),
.B1(net406),
.Y(net397)
);

sky130_fd_sc_hd__mux4_1 c468(
.A0(net130),
.A1(in47),
.A2(net108),
.A3(net259),
.S0(net348),
.S1(net804),
.X(net398)
);

sky130_fd_sc_hd__sdfbbn_1 c469(
.D(net267),
.RESET_B(net395),
.SCD(net404),
.SCE(in13),
.SET_B(net254),
.CLK_N(clk),
.Q(out59),
.Q_N(net399)
);

sky130_fd_sc_hd__a41oi_1 c470(
.A1(net396),
.A2(net410),
.A3(net273),
.A4(net800),
.B1(net807),
.Y(net400)
);

sky130_fd_sc_hd__mux4_4 c471(
.A0(net408),
.A1(out59),
.A2(net410),
.A3(net404),
.S0(net275),
.S1(net755),
.X(net401)
);

sky130_fd_sc_hd__mux4_4 c472(
.A0(net411),
.A1(net393),
.A2(net342),
.A3(net401),
.S0(net399),
.S1(net756),
.X(net402)
);

sky130_fd_sc_hd__mux4_1 c473(
.A0(net412),
.A1(net401),
.A2(net393),
.A3(out41),
.S0(net395),
.S1(net807),
.X(net403)
);

sky130_fd_sc_hd__clkbuf_2 c474(
.A(net788),
.X(out41)
);

sky130_fd_sc_hd__clkinv_1 c475(
.A(net745),
.Y(net404)
);

sky130_fd_sc_hd__clkbuf_1 c476(
.A(net744),
.X(net405)
);

sky130_fd_sc_hd__a21bo_2 c477(
.A1(net19),
.A2(net374),
.B1_N(out53),
.X(net406)
);

sky130_fd_sc_hd__a21boi_0 c478(
.A1(net405),
.A2(net259),
.B1_N(net373),
.Y(net407)
);

sky130_fd_sc_hd__clkinv_16 c479(
.A(net788),
.Y(net408)
);

sky130_fd_sc_hd__clkinv_4 c480(
.A(net788),
.Y(net409)
);

sky130_fd_sc_hd__xor2_1 c481(
.A(net259),
.B(in19),
.X(net410)
);

sky130_fd_sc_hd__dlygate4sd1_1 c482(
.A(net744),
.X(net411)
);

sky130_fd_sc_hd__inv_12 c483(
.A(net747),
.Y(net412)
);

sky130_fd_sc_hd__clkinv_4 c484(
.A(out35),
.Y(out47)
);

sky130_fd_sc_hd__a31oi_4 c485(
.A1(net25),
.A2(out47),
.A3(in39),
.B1(net299),
.Y(net413)
);

sky130_fd_sc_hd__a41o_4 c486(
.A1(in39),
.A2(net307),
.A3(net366),
.A4(out8),
.B1(net299),
.X(net414)
);

sky130_fd_sc_hd__a41o_2 c487(
.A1(net410),
.A2(net308),
.A3(net413),
.A4(net414),
.B1(net799),
.X(net415)
);

sky130_fd_sc_hd__a31o_4 c488(
.A1(net287),
.A2(net415),
.A3(net303),
.B1(net299),
.X(net416)
);

sky130_fd_sc_hd__mux4_4 c489(
.A0(net105),
.A1(net392),
.A2(net303),
.A3(out43),
.S0(net800),
.S1(net807),
.X(net417)
);

sky130_fd_sc_hd__mux2_8 c490(
.A0(net38),
.A1(out45),
.S(net366),
.X(net418)
);

sky130_fd_sc_hd__a41o_4 c491(
.A1(net45),
.A2(net294),
.A3(net418),
.A4(net307),
.B1(net38),
.X(net419)
);

sky130_fd_sc_hd__a41oi_4 c492(
.A1(net351),
.A2(in49),
.A3(out55),
.A4(net268),
.B1(net303),
.Y(net420)
);

sky130_fd_sc_hd__mux4_4 c493(
.A0(net414),
.A1(net418),
.A2(net419),
.A3(out45),
.S0(net417),
.S1(net794),
.X(net421)
);

sky130_fd_sc_hd__buf_12 c494(
.A(out35),
.X(net422)
);

sky130_fd_sc_hd__a41oi_4 c495(
.A1(net308),
.A2(net422),
.A3(out45),
.A4(net410),
.B1(net807),
.Y(net423)
);

sky130_fd_sc_hd__o21ba_1 c496(
.A1(net420),
.A2(net423),
.B1_N(net366),
.X(net424)
);

sky130_fd_sc_hd__o21a_4 c497(
.A1(net303),
.A2(net419),
.B1(net25),
.X(net425)
);

sky130_fd_sc_hd__mux4_2 c498(
.A0(net403),
.A1(net268),
.A2(net423),
.A3(net420),
.S0(net425),
.S1(net807),
.X(net426)
);

sky130_fd_sc_hd__mux4_2 c499(
.A0(net291),
.A1(net105),
.A2(net348),
.A3(in13),
.S0(net425),
.S1(out44),
.X(net427)
);

sky130_fd_sc_hd__mux2_1 c500(
.A0(net424),
.A1(net744),
.S(net809),
.X(net428)
);

sky130_fd_sc_hd__a41oi_1 c501(
.A1(net428),
.A2(net413),
.A3(net414),
.A4(net379),
.B1(net403),
.Y(net429)
);

sky130_fd_sc_hd__a41o_1 c502(
.A1(net423),
.A2(in13),
.A3(net424),
.A4(net425),
.B1(net808),
.X(net430)
);

sky130_fd_sc_hd__o21bai_2 c503(
.A1(net419),
.A2(net424),
.B1_N(net744),
.Y(out25)
);

sky130_fd_sc_hd__a31oi_2 c504(
.A1(net418),
.A2(in39),
.A3(net419),
.B1(net299),
.Y(net431)
);

sky130_fd_sc_hd__clkinv_4 c505(
.A(net742),
.Y(net432)
);

sky130_fd_sc_hd__mux4_2 c526(
.A0(in13),
.A1(out43),
.A2(out54),
.A3(out45),
.S0(out34),
.S1(net796),
.X(out48)
);

sky130_fd_sc_hd__mux4_1 c527(
.A0(net366),
.A1(net294),
.A2(out52),
.A3(out15),
.S0(out48),
.S1(net796),
.X(net433)
);

sky130_fd_sc_hd__xnor2_4 c528(
.A(net209),
.B(net329),
.Y(net434)
);

sky130_fd_sc_hd__clkinv_4 c529(
.A(net731),
.Y(net435)
);

sky130_fd_sc_hd__clkbuf_8 c530(
.A(net731),
.X(net436)
);

sky130_fd_sc_hd__xor2_2 c531(
.A(net201),
.B(net435),
.X(net437)
);

sky130_fd_sc_hd__xnor2_4 c532(
.A(net434),
.B(net435),
.Y(net438)
);

sky130_fd_sc_hd__xnor2_2 c533(
.A(net437),
.B(net435),
.Y(out23)
);

sky130_fd_sc_hd__xnor2_4 c534(
.A(in4),
.B(net81),
.Y(net439)
);

sky130_fd_sc_hd__xor2_2 c535(
.A(net340),
.B(out23),
.X(net440)
);

sky130_fd_sc_hd__a41oi_2 c536(
.A1(net436),
.A2(net332),
.A3(net209),
.A4(net329),
.B1(net218),
.Y(net441)
);

sky130_fd_sc_hd__xor2_2 c537(
.A(net434),
.B(net440),
.X(out39)
);

sky130_fd_sc_hd__xor2_2 c538(
.A(net440),
.B(net771),
.X(net442)
);

sky130_fd_sc_hd__xor2_4 c539(
.A(net438),
.B(out23),
.X(net443)
);

sky130_fd_sc_hd__mux4_1 c540(
.A0(net435),
.A1(net440),
.A2(net340),
.A3(out39),
.S0(net347),
.S1(net802),
.X(net444)
);

sky130_fd_sc_hd__buf_8 c541(
.A(net675),
.X(net445)
);

sky130_fd_sc_hd__a41o_1 c542(
.A1(net329),
.A2(net445),
.A3(net435),
.A4(net443),
.B1(net801),
.X(net446)
);

sky130_fd_sc_hd__inv_12 c543(
.A(net675),
.Y(net447)
);

sky130_fd_sc_hd__a21o_1 c544(
.A1(net439),
.A2(net445),
.B1(out23),
.X(net448)
);

sky130_fd_sc_hd__mux4_2 c545(
.A0(net442),
.A1(net446),
.A2(out39),
.A3(net448),
.S0(net440),
.S1(net434),
.X(net449)
);

sky130_fd_sc_hd__a41oi_2 c546(
.A1(net447),
.A2(net329),
.A3(net332),
.A4(net448),
.B1(net734),
.Y(net450)
);

sky130_fd_sc_hd__buf_8 c547(
.A(net772),
.X(net451)
);

sky130_fd_sc_hd__mux4_2 c548(
.A0(net447),
.A1(net218),
.A2(net340),
.A3(net448),
.S0(net440),
.S1(net442),
.X(net452)
);

sky130_fd_sc_hd__mux4_1 c549(
.A0(net446),
.A1(net448),
.A2(net434),
.A3(in11),
.S0(net734),
.S1(net771),
.X(net453)
);

sky130_fd_sc_hd__o21ai_4 c550(
.A1(net218),
.A2(net448),
.B1(net108),
.Y(net454)
);

sky130_fd_sc_hd__xnor2_4 c551(
.A(net445),
.B(net218),
.Y(net455)
);

sky130_fd_sc_hd__xor2_1 c552(
.A(in11),
.B(net108),
.X(net456)
);

sky130_fd_sc_hd__a31o_2 c553(
.A1(net369),
.A2(net438),
.A3(net79),
.B1(net350),
.X(net457)
);

sky130_fd_sc_hd__xor2_2 c554(
.A(net448),
.B(net353),
.X(net458)
);

sky130_fd_sc_hd__a31oi_1 c555(
.A1(net440),
.A2(net369),
.A3(net446),
.B1(net451),
.Y(net459)
);

sky130_fd_sc_hd__xnor2_2 c556(
.A(net81),
.B(net108),
.Y(net460)
);

sky130_fd_sc_hd__clkinv_16 c557(
.A(net749),
.Y(out24)
);

sky130_fd_sc_hd__a21oi_1 c558(
.A1(net458),
.A2(net460),
.B1(net777),
.Y(net461)
);

sky130_fd_sc_hd__xor2_4 c559(
.A(net772),
.B(net780),
.X(net462)
);

sky130_fd_sc_hd__xnor2_4 c560(
.A(net456),
.B(in0),
.Y(net463)
);

sky130_fd_sc_hd__a21boi_0 c561(
.A1(net463),
.A2(net460),
.B1_N(net780),
.Y(net464)
);

sky130_fd_sc_hd__a41oi_4 c562(
.A1(net357),
.A2(net353),
.A3(net463),
.A4(in0),
.B1(net460),
.Y(net465)
);

sky130_fd_sc_hd__a41oi_2 c563(
.A1(net455),
.A2(net452),
.A3(net464),
.A4(net438),
.B1(net460),
.Y(net466)
);

sky130_fd_sc_hd__a41o_1 c564(
.A1(net465),
.A2(net79),
.A3(out39),
.A4(net218),
.B1(net108),
.X(net467)
);

sky130_fd_sc_hd__o21a_2 c565(
.A1(net463),
.A2(net440),
.B1(net460),
.X(net468)
);

sky130_fd_sc_hd__buf_16 c566(
.A(net749),
.X(net469)
);

sky130_fd_sc_hd__a41o_4 c567(
.A1(net468),
.A2(net334),
.A3(net467),
.A4(net469),
.B1(out8),
.X(net470)
);

sky130_fd_sc_hd__o21ba_1 c568(
.A1(net454),
.A2(net226),
.B1_N(net469),
.X(net471)
);

sky130_fd_sc_hd__clkbuf_2 c569(
.A(net772),
.X(net472)
);

sky130_fd_sc_hd__mux4_1 c570(
.A0(net469),
.A1(net471),
.A2(net357),
.A3(out33),
.S0(in13),
.S1(net746),
.X(net473)
);

sky130_fd_sc_hd__mux4_1 c571(
.A0(net467),
.A1(net369),
.A2(net456),
.A3(in11),
.S0(net469),
.S1(net786),
.X(net474)
);

sky130_fd_sc_hd__a31oi_4 c572(
.A1(net438),
.A2(net748),
.A3(net778),
.B1(net805),
.Y(net475)
);

sky130_fd_sc_hd__a31oi_2 c573(
.A1(net457),
.A2(net70),
.A3(net130),
.B1(net460),
.Y(net476)
);

sky130_fd_sc_hd__o21bai_4 c574(
.A1(net226),
.A2(net469),
.B1_N(net351),
.Y(net477)
);

sky130_fd_sc_hd__a31o_4 c575(
.A1(net70),
.A2(net347),
.A3(net350),
.B1(out22),
.X(net478)
);

sky130_fd_sc_hd__a21o_4 c576(
.A1(net475),
.A2(net347),
.B1(net70),
.X(net479)
);

sky130_fd_sc_hd__o21ai_1 c577(
.A1(net70),
.A2(net748),
.B1(net805),
.Y(net480)
);

sky130_fd_sc_hd__sdfrtp_1 c578(
.D(net390),
.RESET_B(net246),
.SCD(net226),
.SCE(out24),
.CLK(clk),
.Q(net481)
);

sky130_fd_sc_hd__mux4_4 c579(
.A0(net469),
.A1(net481),
.A2(out38),
.A3(net477),
.S0(net478),
.S1(net806),
.X(net482)
);

sky130_fd_sc_hd__sdfbbn_2 c580(
.D(net347),
.RESET_B(in7),
.SCD(net480),
.SCE(net471),
.SET_B(net113),
.CLK_N(clk),
.Q(net484),
.Q_N(net483)
);

sky130_fd_sc_hd__mux4_4 c581(
.A0(net385),
.A1(net347),
.A2(net484),
.A3(net451),
.S0(net457),
.S1(net460),
.X(net485)
);

sky130_fd_sc_hd__clkbuf_16 c582(
.A(net739),
.X(net486)
);

sky130_fd_sc_hd__a41oi_4 c583(
.A1(net486),
.A2(net246),
.A3(net107),
.A4(net350),
.B1(net484),
.Y(net487)
);

sky130_fd_sc_hd__sdfrtp_2 c584(
.D(net477),
.RESET_B(net438),
.SCD(net390),
.SCE(net479),
.CLK(clk),
.Q(net488)
);

sky130_fd_sc_hd__a41oi_1 c585(
.A1(net485),
.A2(net457),
.A3(net488),
.A4(net483),
.B1(net469),
.Y(net489)
);

sky130_fd_sc_hd__a41oi_4 c586(
.A1(net446),
.A2(net462),
.A3(net70),
.A4(net460),
.B1(net477),
.Y(net490)
);

sky130_fd_sc_hd__a41o_1 c587(
.A1(net480),
.A2(net481),
.A3(net484),
.A4(net347),
.B1(out30),
.X(net491)
);

sky130_fd_sc_hd__mux4_4 c588(
.A0(net487),
.A1(net477),
.A2(net351),
.A3(net130),
.S0(net469),
.S1(net471),
.X(net492)
);

sky130_fd_sc_hd__sdfrtp_4 c589(
.D(net452),
.RESET_B(net385),
.SCD(net488),
.SCE(out30),
.CLK(clk),
.Q(net493)
);

sky130_fd_sc_hd__a41oi_2 c590(
.A1(net477),
.A2(net493),
.A3(net1),
.A4(net488),
.B1(out22),
.Y(net494)
);

sky130_fd_sc_hd__a31o_1 c591(
.A1(net491),
.A2(net494),
.A3(net70),
.B1(net130),
.X(net495)
);

sky130_fd_sc_hd__a41oi_2 c592(
.A1(net462),
.A2(net493),
.A3(net481),
.A4(net483),
.B1(net778),
.Y(net496)
);

sky130_fd_sc_hd__mux4_4 c593(
.A0(net496),
.A1(net347),
.A2(net451),
.A3(out7),
.S0(net493),
.S1(net731),
.X(net497)
);

sky130_fd_sc_hd__a31o_1 c594(
.A1(net270),
.A2(net351),
.A3(net488),
.B1(net777),
.X(net498)
);

sky130_fd_sc_hd__a31oi_4 c595(
.A1(net481),
.A2(out33),
.A3(out39),
.B1(net483),
.Y(net499)
);

sky130_fd_sc_hd__a31oi_4 c596(
.A1(net482),
.A2(net391),
.A3(out39),
.B1(net777),
.Y(net500)
);

sky130_fd_sc_hd__o21bai_1 c597(
.A1(net105),
.A2(net404),
.B1_N(net756),
.Y(net501)
);

sky130_fd_sc_hd__sdfbbp_1 c598(
.D(net500),
.RESET_B(net501),
.SCD(net494),
.SCE(net452),
.SET_B(net391),
.CLK(clk),
.Q(out0),
.Q_N(net502)
);

sky130_fd_sc_hd__a31oi_4 c599(
.A1(net493),
.A2(net1),
.A3(out24),
.B1(net501),
.Y(net503)
);

sky130_fd_sc_hd__a41oi_2 c600(
.A1(out41),
.A2(net1),
.A3(net493),
.A4(net460),
.B1(net806),
.Y(net504)
);

sky130_fd_sc_hd__a31o_1 c601(
.A1(net1),
.A2(net504),
.A3(out38),
.B1(net502),
.X(net505)
);

sky130_fd_sc_hd__mux4_1 c602(
.A0(net500),
.A1(net505),
.A2(out0),
.A3(out38),
.S0(net494),
.S1(net748),
.X(net506)
);

sky130_fd_sc_hd__o21bai_4 c603(
.A1(net504),
.A2(net402),
.B1_N(out24),
.Y(net507)
);

sky130_fd_sc_hd__mux4_2 c604(
.A0(net498),
.A1(net493),
.A2(net501),
.A3(net497),
.S0(out23),
.S1(net782),
.X(net508)
);

sky130_fd_sc_hd__clkinv_1 c605(
.A(net743),
.Y(net509)
);

sky130_fd_sc_hd__a31oi_2 c606(
.A1(out24),
.A2(net481),
.A3(net768),
.B1(net782),
.Y(net510)
);

sky130_fd_sc_hd__inv_8 c607(
.A(net743),
.Y(out31)
);

sky130_fd_sc_hd__mux2_8 c608(
.A0(net451),
.A1(net501),
.S(net494),
.X(net511)
);

sky130_fd_sc_hd__sdfbbn_1 c609(
.D(net488),
.RESET_B(net497),
.SCD(net501),
.SCE(net511),
.SET_B(net507),
.CLK_N(clk),
.Q(net513),
.Q_N(net512)
);

sky130_fd_sc_hd__sdfbbn_2 c610(
.D(net503),
.RESET_B(out0),
.SCD(net511),
.SCE(net512),
.SET_B(net460),
.CLK_N(clk),
.Q(net515),
.Q_N(net514)
);

sky130_fd_sc_hd__a31o_1 c611(
.A1(net509),
.A2(net379),
.A3(net515),
.B1(in33),
.X(net516)
);

sky130_fd_sc_hd__mux4_2 c612(
.A0(net515),
.A1(in7),
.A2(out24),
.A3(net404),
.S0(net452),
.S1(net108),
.X(net517)
);

sky130_fd_sc_hd__mux4_2 c613(
.A0(net501),
.A1(net514),
.A2(net12),
.A3(net395),
.S0(net512),
.S1(net782),
.X(net518)
);

sky130_fd_sc_hd__a41oi_4 c614(
.A1(net518),
.A2(net460),
.A3(net512),
.A4(out23),
.B1(net777),
.Y(net519)
);

sky130_fd_sc_hd__mux4_4 c615(
.A0(net511),
.A1(out26),
.A2(net518),
.A3(net504),
.S0(net756),
.S1(net777),
.X(net520)
);

sky130_fd_sc_hd__sdfbbp_1 c616(
.D(net395),
.RESET_B(net513),
.SCD(net12),
.SCE(net478),
.SET_B(net518),
.CLK(clk),
.Q(net522),
.Q_N(net521)
);

sky130_fd_sc_hd__mux4_2 c617(
.A0(out37),
.A1(net509),
.A2(net521),
.A3(net425),
.S0(net452),
.S1(net809),
.X(net523)
);

sky130_fd_sc_hd__mux4_1 c618(
.A0(net404),
.A1(net12),
.A2(net161),
.A3(out37),
.S0(in33),
.S1(in13),
.X(net524)
);

sky130_fd_sc_hd__mux4_4 c619(
.A0(net510),
.A1(out8),
.A2(net391),
.A3(out37),
.S0(net404),
.S1(net778),
.X(net525)
);

sky130_fd_sc_hd__mux4_1 c620(
.A0(net522),
.A1(net460),
.A2(net417),
.A3(net425),
.S0(out37),
.S1(net161),
.X(net526)
);

sky130_fd_sc_hd__a41o_1 c621(
.A1(net417),
.A2(out15),
.A3(out38),
.A4(out18),
.B1(out37),
.X(net527)
);

sky130_fd_sc_hd__mux4_2 c622(
.A0(net161),
.A1(net480),
.A2(net12),
.A3(net513),
.S0(in49),
.S1(out21),
.X(net528)
);

sky130_fd_sc_hd__mux4_4 c623(
.A0(out26),
.A1(net522),
.A2(net264),
.A3(out39),
.S0(in49),
.S1(net768),
.X(net529)
);

sky130_fd_sc_hd__mux4_4 c624(
.A0(net518),
.A1(out18),
.A2(out26),
.A3(net513),
.S0(net521),
.S1(in49),
.X(net530)
);

sky130_fd_sc_hd__a41oi_2 c625(
.A1(net480),
.A2(net12),
.A3(net529),
.A4(out18),
.B1(net522),
.Y(net531)
);

sky130_fd_sc_hd__mux4_2 c626(
.A0(net525),
.A1(net478),
.A2(net379),
.A3(net518),
.S0(net521),
.S1(out31),
.X(net532)
);

sky130_fd_sc_hd__mux4_1 c627(
.A0(net422),
.A1(out37),
.A2(net478),
.A3(net514),
.S0(net809),
.S1(net811),
.X(net533)
);

sky130_fd_sc_hd__mux4_2 c628(
.A0(net422),
.A1(out37),
.A2(net478),
.A3(net768),
.S0(out2),
.S1(net811),
.X(out32)
);

sky130_fd_sc_hd__mux4_2 c629(
.A0(net392),
.A1(out24),
.A2(out23),
.A3(out7),
.S0(in33),
.S1(net760),
.X(net534)
);

sky130_fd_sc_hd__mux4_4 c630(
.A0(net529),
.A1(net509),
.A2(in49),
.A3(net513),
.S0(net268),
.S1(net478),
.X(net535)
);

sky130_fd_sc_hd__mux4_4 c631(
.A0(net528),
.A1(net533),
.A2(net522),
.A3(out26),
.S0(net514),
.S1(net811),
.X(out29)
);

sky130_fd_sc_hd__mux4_1 c632(
.A0(in49),
.A1(out32),
.A2(net480),
.A3(net105),
.S0(net761),
.S1(net778),
.X(net536)
);

sky130_fd_sc_hd__mux4_1 c633(
.A0(net379),
.A1(net392),
.A2(net533),
.A3(net169),
.S0(out37),
.S1(net811),
.X(net537)
);

sky130_fd_sc_hd__a41oi_1 c634(
.A1(net478),
.A2(out32),
.A3(out37),
.A4(net395),
.B1(net525),
.Y(net538)
);

sky130_fd_sc_hd__mux4_4 c635(
.A0(net536),
.A1(net515),
.A2(net538),
.A3(out15),
.S0(net379),
.S1(net812),
.X(net539)
);

sky130_fd_sc_hd__mux4_4 c636(
.A0(net534),
.A1(out32),
.A2(net478),
.A3(out37),
.S0(net811),
.S1(net812),
.X(net540)
);

sky130_fd_sc_hd__mux4_2 c637(
.A0(net524),
.A1(net540),
.A2(net538),
.A3(net533),
.S0(net778),
.S1(out21),
.X(net541)
);

sky130_fd_sc_hd__o21ba_1 c660(
.A1(net217),
.A2(net207),
.B1_N(net435),
.X(net542)
);

sky130_fd_sc_hd__a21bo_2 c661(
.A1(net218),
.A2(net69),
.B1_N(net330),
.X(net543)
);

sky130_fd_sc_hd__o21ai_4 c662(
.A1(net211),
.A2(in14),
.B1(net435),
.Y(net544)
);

sky130_fd_sc_hd__clkinv_4 c663(
.A(net746),
.Y(net545)
);

sky130_fd_sc_hd__xnor2_2 c664(
.A(net77),
.B(net435),
.Y(net546)
);

sky130_fd_sc_hd__xnor2_1 c665(
.A(in14),
.B(net69),
.Y(net547)
);

sky130_fd_sc_hd__a21o_4 c666(
.A1(net69),
.A2(net77),
.B1(net435),
.X(net548)
);

sky130_fd_sc_hd__xnor2_2 c667(
.A(net435),
.B(net69),
.Y(net549)
);

sky130_fd_sc_hd__xnor2_4 c668(
.A(net547),
.B(net545),
.Y(net550)
);

sky130_fd_sc_hd__xnor2_4 c669(
.A(net550),
.B(net547),
.Y(net551)
);

sky130_fd_sc_hd__xor2_1 c670(
.A(net545),
.B(net551),
.X(net552)
);

sky130_fd_sc_hd__o21ai_4 c671(
.A1(net326),
.A2(net547),
.B1(net546),
.Y(net553)
);

sky130_fd_sc_hd__mux4_4 c672(
.A0(net207),
.A1(net551),
.A2(net553),
.A3(in14),
.S0(net550),
.S1(net452),
.X(net554)
);

sky130_fd_sc_hd__xor2_2 c673(
.A(net211),
.B(net553),
.X(net555)
);

sky130_fd_sc_hd__dlygate4sd1_1 c674(
.A(net746),
.X(net556)
);

sky130_fd_sc_hd__mux4_2 c675(
.A0(net552),
.A1(net556),
.A2(net544),
.A3(net543),
.S0(net549),
.S1(net435),
.X(net557)
);

sky130_fd_sc_hd__xnor2_2 c676(
.A(net326),
.B(out21),
.Y(net558)
);

sky130_fd_sc_hd__o21bai_1 c677(
.A1(net555),
.A2(net549),
.B1_N(net553),
.Y(net559)
);

sky130_fd_sc_hd__mux4_1 c678(
.A0(net555),
.A1(net558),
.A2(net543),
.A3(net556),
.S0(net334),
.S1(net553),
.X(net560)
);

sky130_fd_sc_hd__a41oi_4 c679(
.A1(net558),
.A2(net556),
.A3(net546),
.A4(in14),
.B1(net784),
.Y(net561)
);

sky130_fd_sc_hd__mux4_4 c680(
.A0(net549),
.A1(net545),
.A2(net552),
.A3(net207),
.S0(net555),
.S1(net784),
.X(net562)
);

sky130_fd_sc_hd__mux4_4 c681(
.A0(net561),
.A1(net562),
.A2(net452),
.A3(net556),
.S0(net334),
.S1(net784),
.X(net563)
);

sky130_fd_sc_hd__sdfsbp_1 c682(
.D(net556),
.SCD(net334),
.SCE(net551),
.SET_B(net559),
.CLK(clk),
.Q(net565),
.Q_N(net564)
);

sky130_fd_sc_hd__o21bai_1 c683(
.A1(net472),
.A2(in13),
.B1_N(net105),
.Y(net566)
);

sky130_fd_sc_hd__o21a_1 c684(
.A1(net553),
.A2(out21),
.B1(net802),
.X(net567)
);

sky130_fd_sc_hd__a21oi_2 c685(
.A1(net565),
.A2(in33),
.B1(net542),
.Y(net568)
);

sky130_fd_sc_hd__sdfsbp_2 c686(
.D(net107),
.SCD(net568),
.SCE(net471),
.SET_B(net558),
.CLK(clk),
.Q(net570),
.Q_N(net569)
);

sky130_fd_sc_hd__xnor2_2 c687(
.A(net570),
.B(net542),
.Y(net571)
);

sky130_fd_sc_hd__a21bo_2 c688(
.A1(net546),
.A2(net571),
.B1_N(net350),
.X(net572)
);

sky130_fd_sc_hd__mux4_1 c689(
.A0(net549),
.A1(net570),
.A2(net452),
.A3(net571),
.S0(net551),
.S1(net330),
.X(net573)
);

sky130_fd_sc_hd__mux2_8 c690(
.A0(net567),
.A1(net569),
.S(net786),
.X(net574)
);

sky130_fd_sc_hd__a21bo_2 c691(
.A1(net564),
.A2(net556),
.B1_N(out21),
.X(net575)
);

sky130_fd_sc_hd__a41oi_4 c692(
.A1(net334),
.A2(net570),
.A3(net471),
.A4(net452),
.B1(net218),
.Y(net576)
);

sky130_fd_sc_hd__a21o_4 c693(
.A1(net542),
.A2(net571),
.B1(net574),
.X(net577)
);

sky130_fd_sc_hd__clkbuf_4 c694(
.A(net766),
.X(net578)
);

sky130_fd_sc_hd__inv_8 c695(
.A(net766),
.Y(net579)
);

sky130_fd_sc_hd__mux4_2 c696(
.A0(net567),
.A1(net575),
.A2(net579),
.A3(net472),
.S0(net548),
.S1(net718),
.X(net580)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c697(
.A(net779),
.X(net581)
);

sky130_fd_sc_hd__mux4_4 c698(
.A0(net577),
.A1(net351),
.A2(net334),
.A3(net544),
.S0(net464),
.S1(net575),
.X(net582)
);

sky130_fd_sc_hd__a21bo_1 c699(
.A1(net464),
.A2(net581),
.B1_N(net571),
.X(net583)
);

sky130_fd_sc_hd__a41oi_1 c700(
.A1(net579),
.A2(net583),
.A3(net464),
.A4(out8),
.B1(net770),
.Y(net584)
);

sky130_fd_sc_hd__a41o_1 c701(
.A1(net580),
.A2(net569),
.A3(net577),
.A4(net564),
.B1(net784),
.X(net585)
);

sky130_fd_sc_hd__mux4_4 c702(
.A0(net566),
.A1(net461),
.A2(net579),
.A3(net571),
.S0(net770),
.S1(net784),
.X(net586)
);

sky130_fd_sc_hd__a41oi_1 c703(
.A1(net549),
.A2(net575),
.A3(net718),
.A4(net784),
.B1(net814),
.Y(out4)
);

sky130_fd_sc_hd__a31o_4 c704(
.A1(net574),
.A2(net330),
.A3(net484),
.B1(net814),
.X(net587)
);

sky130_fd_sc_hd__a41o_2 c705(
.A1(net548),
.A2(net544),
.A3(net373),
.A4(net484),
.B1(net587),
.X(net588)
);

sky130_fd_sc_hd__mux4_1 c706(
.A0(out7),
.A1(net452),
.A2(net107),
.A3(net548),
.S0(net805),
.S1(net814),
.X(net589)
);

sky130_fd_sc_hd__sdfbbn_1 c707(
.D(net578),
.RESET_B(net373),
.SCD(net130),
.SCE(in7),
.SET_B(net815),
.CLK_N(clk),
.Q(net591),
.Q_N(net590)
);

sky130_fd_sc_hd__a41oi_4 c708(
.A1(net559),
.A2(net547),
.A3(net581),
.A4(net113),
.B1(net787),
.Y(net592)
);

sky130_fd_sc_hd__sdfbbn_2 c709(
.D(net553),
.RESET_B(net471),
.SCD(net460),
.SCE(net330),
.SET_B(out16),
.CLK_N(clk),
.Q(net594),
.Q_N(net593)
);

sky130_fd_sc_hd__a41o_1 c710(
.A1(net594),
.A2(net0),
.A3(out4),
.A4(net574),
.B1(net483),
.X(net595)
);

sky130_fd_sc_hd__a31o_1 c711(
.A1(net595),
.A2(net594),
.A3(net553),
.B1(net813),
.X(net596)
);

sky130_fd_sc_hd__a41oi_2 c712(
.A1(net351),
.A2(net551),
.A3(net479),
.A4(net735),
.B1(net814),
.Y(net597)
);

sky130_fd_sc_hd__mux4_1 c713(
.A0(net587),
.A1(net591),
.A2(net483),
.A3(net593),
.S0(net787),
.S1(net815),
.X(net598)
);

sky130_fd_sc_hd__mux4_4 c714(
.A0(net578),
.A1(net594),
.A2(in7),
.A3(net735),
.S0(out19),
.S1(net787),
.X(net599)
);

sky130_fd_sc_hd__mux4_4 c715(
.A0(net599),
.A1(net330),
.A2(net460),
.A3(net814),
.S0(net815),
.S1(net816),
.X(net600)
);

sky130_fd_sc_hd__a41oi_1 c716(
.A1(net600),
.A2(net547),
.A3(net108),
.A4(net593),
.B1(net596),
.Y(net601)
);

sky130_fd_sc_hd__a41oi_2 c717(
.A1(net2),
.A2(net594),
.A3(net330),
.A4(net590),
.B1(net548),
.Y(net602)
);

sky130_fd_sc_hd__a41oi_4 c718(
.A1(net596),
.A2(net593),
.A3(net787),
.A4(net805),
.B1(net816),
.Y(net603)
);

sky130_fd_sc_hd__mux4_2 c719(
.A0(net455),
.A1(net594),
.A2(net603),
.A3(net544),
.S0(out19),
.S1(net786),
.X(net604)
);

sky130_fd_sc_hd__mux4_4 c720(
.A0(net604),
.A1(net596),
.A2(net559),
.A3(net484),
.S0(net581),
.S1(net108),
.X(net605)
);

sky130_fd_sc_hd__mux4_4 c721(
.A0(net596),
.A1(net2),
.A2(net604),
.A3(net593),
.S0(net483),
.S1(net818),
.X(net606)
);

sky130_fd_sc_hd__mux4_2 c722(
.A0(net471),
.A1(net583),
.A2(net604),
.A3(net590),
.S0(net818),
.S1(net819),
.X(net607)
);

sky130_fd_sc_hd__mux4_1 c723(
.A0(net604),
.A1(net330),
.A2(net816),
.A3(net818),
.S0(net820),
.S1(net822),
.X(net608)
);

sky130_fd_sc_hd__mux4_1 c724(
.A0(net551),
.A1(net600),
.A2(net604),
.A3(net817),
.S0(net819),
.S1(net822),
.X(net609)
);

sky130_fd_sc_hd__mux4_1 c725(
.A0(net574),
.A1(net565),
.A2(net604),
.A3(net733),
.S0(net817),
.S1(net821),
.X(net610)
);

sky130_fd_sc_hd__a31o_2 c726(
.A1(net479),
.A2(net460),
.A3(net568),
.B1(net397),
.X(net611)
);

sky130_fd_sc_hd__mux4_1 c727(
.A0(net0),
.A1(net568),
.A2(net544),
.A3(net590),
.S0(net780),
.S1(net823),
.X(net612)
);

sky130_fd_sc_hd__mux2_4 c728(
.A0(net0),
.A1(out0),
.S(net779),
.X(net613)
);

sky130_fd_sc_hd__mux4_4 c729(
.A0(net373),
.A1(net591),
.A2(net452),
.A3(net780),
.S0(net813),
.S1(net816),
.X(net614)
);

sky130_fd_sc_hd__mux4_2 c730(
.A0(net484),
.A1(net452),
.A2(net558),
.A3(out16),
.S0(net810),
.S1(net813),
.X(net615)
);

sky130_fd_sc_hd__sdfstp_1 c731(
.D(net612),
.SCD(net479),
.SCE(net452),
.SET_B(out9),
.CLK(clk),
.Q(net616)
);

sky130_fd_sc_hd__a41o_2 c732(
.A1(net544),
.A2(out4),
.A3(net2),
.A4(out0),
.B1(net815),
.X(out10)
);

sky130_fd_sc_hd__o21bai_4 c733(
.A1(net494),
.A2(net813),
.B1_N(net823),
.Y(net617)
);

sky130_fd_sc_hd__mux4_4 c734(
.A0(net394),
.A1(net617),
.A2(net351),
.A3(net397),
.S0(net616),
.S1(net816),
.X(net618)
);

sky130_fd_sc_hd__mux4_1 c735(
.A0(net460),
.A1(net108),
.A2(out4),
.A3(out10),
.S0(net816),
.S1(net823),
.X(net619)
);

sky130_fd_sc_hd__a41oi_2 c736(
.A1(net130),
.A2(net617),
.A3(net479),
.A4(net733),
.B1(net824),
.Y(net620)
);

sky130_fd_sc_hd__sdfbbp_1 c737(
.D(net602),
.RESET_B(net617),
.SCD(net568),
.SCE(net373),
.SET_B(in33),
.CLK(clk),
.Q(net622),
.Q_N(net621)
);

sky130_fd_sc_hd__a41oi_4 c738(
.A1(net596),
.A2(net616),
.A3(net621),
.A4(out10),
.B1(net568),
.Y(net623)
);

sky130_fd_sc_hd__mux4_1 c739(
.A0(net622),
.A1(net113),
.A2(net397),
.A3(net616),
.S0(net780),
.S1(net824),
.X(net624)
);

sky130_fd_sc_hd__mux4_2 c740(
.A0(out4),
.A1(net616),
.A2(net558),
.A3(net779),
.S0(net813),
.S1(net816),
.X(net625)
);

sky130_fd_sc_hd__mux4_2 c741(
.A0(net617),
.A1(net581),
.A2(net568),
.A3(net616),
.S0(out10),
.S1(net813),
.X(net626)
);

sky130_fd_sc_hd__mux4_4 c742(
.A0(net625),
.A1(net558),
.A2(net394),
.A3(out16),
.S0(net776),
.S1(net785),
.X(out12)
);

sky130_fd_sc_hd__mux4_1 c743(
.A0(net624),
.A1(net616),
.A2(out18),
.A3(net785),
.S0(net821),
.S1(net824),
.X(net627)
);

sky130_fd_sc_hd__a41oi_2 c744(
.A1(net616),
.A2(net479),
.A3(net731),
.A4(net776),
.B1(net824),
.Y(net628)
);

sky130_fd_sc_hd__a41oi_2 c745(
.A1(net603),
.A2(net108),
.A3(net544),
.A4(net621),
.B1(net766),
.Y(net629)
);

sky130_fd_sc_hd__a31o_2 c746(
.A1(net113),
.A2(net351),
.A3(net766),
.B1(net824),
.X(net630)
);

sky130_fd_sc_hd__mux4_1 c747(
.A0(net629),
.A1(out59),
.A2(net602),
.A3(out12),
.S0(net373),
.S1(net616),
.X(net631)
);

sky130_fd_sc_hd__mux4_2 c748(
.A0(net613),
.A1(net538),
.A2(net113),
.A3(net460),
.S0(out10),
.S1(out2),
.X(net632)
);

sky130_fd_sc_hd__mux4_2 c749(
.A0(net591),
.A1(net558),
.A2(out7),
.A3(in33),
.S0(net350),
.S1(net811),
.X(net633)
);

sky130_fd_sc_hd__a41o_1 c750(
.A1(net113),
.A2(net558),
.A3(net538),
.A4(out17),
.B1(net815),
.X(net634)
);

sky130_fd_sc_hd__mux4_4 c751(
.A0(net558),
.A1(out18),
.A2(net581),
.A3(net460),
.S0(out10),
.S1(net822),
.X(net635)
);

sky130_fd_sc_hd__mux4_4 c752(
.A0(net452),
.A1(out59),
.A2(net558),
.A3(out7),
.S0(net775),
.S1(net811),
.X(net636)
);

sky130_fd_sc_hd__mux4_4 c753(
.A0(net633),
.A1(net415),
.A2(net397),
.A3(out10),
.S0(net776),
.S1(net810),
.X(net637)
);

sky130_fd_sc_hd__mux4_2 c754(
.A0(net425),
.A1(net158),
.A2(net432),
.A3(out10),
.S0(net460),
.S1(net812),
.X(net638)
);

sky130_fd_sc_hd__mux4_4 c755(
.A0(net633),
.A1(out8),
.A2(net415),
.A3(net399),
.S0(out5),
.S1(net769),
.X(net639)
);

sky130_fd_sc_hd__mux4_1 c756(
.A0(net105),
.A1(net633),
.A2(net502),
.A3(net397),
.S0(net538),
.S1(net820),
.X(net640)
);

sky130_fd_sc_hd__mux4_4 c757(
.A0(net432),
.A1(out59),
.A2(net105),
.A3(out5),
.S0(out17),
.S1(net815),
.X(net641)
);

sky130_fd_sc_hd__mux4_2 c758(
.A0(net415),
.A1(net581),
.A2(out15),
.A3(net785),
.S0(net810),
.S1(net823),
.X(net642)
);

sky130_fd_sc_hd__mux4_4 c759(
.A0(out7),
.A1(net633),
.A2(net460),
.A3(net397),
.S0(net761),
.S1(out1),
.X(net643)
);

sky130_fd_sc_hd__mux4_4 c760(
.A0(out8),
.A1(in33),
.A2(net775),
.A3(net785),
.S0(net812),
.S1(net823),
.X(net644)
);

sky130_fd_sc_hd__mux4_4 c761(
.A0(net158),
.A1(net622),
.A2(net633),
.A3(net399),
.S0(net452),
.S1(out2),
.X(net645)
);

sky130_fd_sc_hd__mux4_4 c762(
.A0(net169),
.A1(out12),
.A2(net425),
.A3(net769),
.S0(net823),
.S1(net825),
.X(net646)
);

sky130_fd_sc_hd__mux4_4 c763(
.A0(net397),
.A1(in33),
.A2(out15),
.A3(net776),
.S0(net785),
.S1(net825),
.X(net647)
);

sky130_fd_sc_hd__mux4_1 c764(
.A0(net397),
.A1(net644),
.A2(net432),
.A3(net425),
.S0(net558),
.S1(net825),
.X(net648)
);

sky130_fd_sc_hd__mux4_2 c765(
.A0(net630),
.A1(net641),
.A2(net351),
.A3(net502),
.S0(out9),
.S1(out3),
.X(net649)
);

sky130_fd_sc_hd__mux4_1 c766(
.A0(net419),
.A1(net432),
.A2(out10),
.A3(net815),
.S0(net825),
.S1(out3),
.X(net650)
);

sky130_fd_sc_hd__mux4_2 c767(
.A0(net643),
.A1(net649),
.A2(out10),
.A3(out4),
.S0(net399),
.S1(out3),
.X(net651)
);

sky130_fd_sc_hd__mux4_1 c768(
.A0(net397),
.A1(net643),
.A2(out11),
.A3(out5),
.S0(net825),
.S1(out3),
.X(net652)
);

sky130_fd_sc_hd__mux4_4 c769(
.A0(net452),
.A1(net415),
.A2(net502),
.A3(out30),
.S0(out19),
.S1(net785),
.X(net653)
);

sky130_fd_sc_hd__a41oi_2 merge790(
.A1(net163),
.A2(net68),
.A3(out45),
.A4(net6),
.B1(net311),
.Y(net654)
);

sky130_fd_sc_hd__mux4_4 merge791(
.A0(net182),
.A1(net29),
.A2(net52),
.A3(net167),
.S0(net139),
.S1(out15),
.X(net655)
);

sky130_fd_sc_hd__a41oi_1 merge792(
.A1(net272),
.A2(net273),
.A3(net274),
.A4(net254),
.B1(net268),
.Y(net656)
);

sky130_fd_sc_hd__a41o_2 merge793(
.A1(net543),
.A2(net435),
.A3(net219),
.A4(net552),
.B1(net452),
.X(net657)
);

sky130_fd_sc_hd__mux4_4 merge794(
.A0(net116),
.A1(net115),
.A2(net3),
.A3(net131),
.S0(net125),
.S1(out15),
.X(net658)
);

sky130_fd_sc_hd__a41o_2 merge795(
.A1(net571),
.A2(net577),
.A3(net569),
.A4(net572),
.B1(in13),
.X(net659)
);

sky130_fd_sc_hd__mux4_2 merge796(
.A0(net330),
.A1(net452),
.A2(in0),
.A3(net467),
.S0(net746),
.S1(net801),
.X(net660)
);

sky130_fd_sc_hd__a31o_2 merge797(
.A1(net332),
.A2(net326),
.A3(net327),
.B1(net334),
.X(net661)
);

sky130_fd_sc_hd__mux4_1 merge798(
.A0(net348),
.A1(net403),
.A2(net421),
.A3(net105),
.S0(net303),
.S1(net794),
.X(net662)
);

sky130_fd_sc_hd__a31oi_4 merge799(
.A1(net243),
.A2(out18),
.A3(net247),
.B1(net254),
.Y(net663)
);

sky130_fd_sc_hd__mux4_2 merge800(
.A0(net507),
.A1(out15),
.A2(net508),
.A3(net505),
.S0(net479),
.S1(net768),
.X(net664)
);

sky130_fd_sc_hd__a41o_2 merge801(
.A1(net254),
.A2(net406),
.A3(net155),
.A4(net19),
.B1(net806),
.X(net665)
);

sky130_fd_sc_hd__a31oi_1 merge802(
.A1(net56),
.A2(in45),
.A3(net55),
.B1(net791),
.Y(net666)
);

sky130_fd_sc_hd__a31oi_1 merge803(
.A1(net170),
.A2(net25),
.A3(net166),
.B1(net737),
.Y(net667)
);

sky130_fd_sc_hd__a41o_1 merge804(
.A1(net223),
.A2(net224),
.A3(net214),
.A4(net228),
.B1(net83),
.X(net668)
);

sky130_fd_sc_hd__a41o_4 merge805(
.A1(net331),
.A2(net228),
.A3(net205),
.A4(net92),
.B1(net695),
.X(net669)
);

sky130_fd_sc_hd__a41o_2 merge806(
.A1(net90),
.A2(net213),
.A3(net217),
.A4(net219),
.B1(net797),
.X(net670)
);

sky130_fd_sc_hd__a31oi_2 merge807(
.A1(net228),
.A2(net259),
.A3(net372),
.B1(out15),
.Y(net671)
);

sky130_fd_sc_hd__a31oi_1 merge808(
.A1(net332),
.A2(net86),
.A3(net334),
.B1(net801),
.Y(net672)
);

sky130_fd_sc_hd__a31o_1 merge809(
.A1(net384),
.A2(net379),
.A3(net256),
.B1(net247),
.X(net673)
);

sky130_fd_sc_hd__mux4_1 merge810(
.A0(net188),
.A1(net179),
.A2(net49),
.A3(net296),
.S0(net302),
.S1(net299),
.X(net674)
);

sky130_fd_sc_hd__buf_8 merge811(
.A(net747),
.X(net675)
);

sky130_fd_sc_hd__mux4_4 merge812(
.A0(net359),
.A1(net92),
.A2(net350),
.A3(net452),
.S0(out18),
.S1(net778),
.X(net676)
);

sky130_fd_sc_hd__mux4_1 merge813(
.A0(net464),
.A1(net471),
.A2(net445),
.A3(net86),
.S0(net444),
.S1(net780),
.X(net677)
);

sky130_fd_sc_hd__mux4_2 merge814(
.A0(net3),
.A1(net130),
.A2(net114),
.A3(net236),
.S0(out33),
.S1(net107),
.X(net678)
);

sky130_fd_sc_hd__mux4_4 merge815(
.A0(in47),
.A1(net254),
.A2(net12),
.A3(net311),
.S0(net68),
.S1(net763),
.X(net679)
);

sky130_fd_sc_hd__mux4_1 merge816(
.A0(net146),
.A1(net152),
.A2(net7),
.A3(net182),
.S0(net186),
.S1(net722),
.X(net680)
);

sky130_fd_sc_hd__mux4_2 merge817(
.A0(net374),
.A1(net25),
.A2(net254),
.A3(net315),
.S0(net199),
.S1(net293),
.X(net681)
);

sky130_fd_sc_hd__a41o_4 merge818(
.A1(net267),
.A2(net273),
.A3(net264),
.A4(net755),
.B1(net806),
.X(net682)
);

sky130_fd_sc_hd__mux4_1 merge819(
.A0(net56),
.A1(net52),
.A2(net185),
.A3(net68),
.S0(net167),
.S1(net789),
.X(net683)
);

sky130_fd_sc_hd__mux4_2 merge820(
.A0(net245),
.A1(net123),
.A2(net130),
.A3(net431),
.S0(out25),
.S1(net808),
.X(net684)
);

sky130_fd_sc_hd__a41o_4 merge821(
.A1(in19),
.A2(net201),
.A3(net325),
.A4(net346),
.B1(net343),
.X(net685)
);

sky130_fd_sc_hd__mux4_1 merge822(
.A0(net348),
.A1(net107),
.A2(net362),
.A3(net409),
.S0(out41),
.S1(net273),
.X(net686)
);

sky130_fd_sc_hd__mux4_1 merge823(
.A0(net461),
.A1(net579),
.A2(net105),
.A3(net343),
.S0(net358),
.S1(net362),
.X(net687)
);

sky130_fd_sc_hd__mux4_1 merge824(
.A0(net93),
.A1(net368),
.A2(net364),
.A3(net443),
.S0(net444),
.S1(net446),
.X(net688)
);

sky130_fd_sc_hd__xor2_4 merge825(
.A(net614),
.B(net615),
.X(net689)
);

sky130_fd_sc_hd__xnor2_4 merge826(
.A(net426),
.B(net429),
.Y(net690)
);

sky130_fd_sc_hd__xor2_4 merge827(
.A(net149),
.B(net680),
.X(net691)
);

sky130_fd_sc_hd__xor2_1 merge828(
.A(net288),
.B(net298),
.X(net692)
);

sky130_fd_sc_hd__xor2_2 merge829(
.A(net517),
.B(net519),
.X(net693)
);

sky130_fd_sc_hd__dfrbp_1 merge830(
.D(net337),
.RESET_B(net661),
.CLK(clk),
.Q(net695),
.Q_N(net694)
);

sky130_fd_sc_hd__xor2_1 merge831(
.A(net164),
.B(net667),
.X(net696)
);

sky130_fd_sc_hd__dfrbp_2 merge832(
.D(net187),
.RESET_B(net655),
.CLK(clk),
.Q(out49),
.Q_N(net697)
);

sky130_fd_sc_hd__xnor2_1 merge833(
.A(net470),
.B(net459),
.Y(net698)
);

sky130_fd_sc_hd__xnor2_1 merge834(
.A(net554),
.B(net557),
.Y(net699)
);

sky130_fd_sc_hd__xnor2_2 merge835(
.A(net526),
.B(net530),
.Y(net700)
);

sky130_fd_sc_hd__xor2_1 merge836(
.A(net237),
.B(net230),
.X(net701)
);

sky130_fd_sc_hd__xor2_2 merge837(
.A(net449),
.B(net450),
.X(net702)
);

sky130_fd_sc_hd__dfrtn_1 merge838(
.D(net670),
.RESET_B(net216),
.CLK_N(clk),
.Q(net703)
);

sky130_fd_sc_hd__dfrtp_1 merge839(
.D(net588),
.RESET_B(net592),
.CLK(clk),
.Q(out16)
);

sky130_fd_sc_hd__xnor2_2 merge840(
.A(net489),
.B(net490),
.Y(net704)
);

sky130_fd_sc_hd__xor2_4 merge841(
.A(net354),
.B(net370),
.X(net705)
);

sky130_fd_sc_hd__xor2_1 merge842(
.A(net381),
.B(net380),
.X(net706)
);

sky130_fd_sc_hd__xor2_4 merge843(
.A(net666),
.B(net683),
.X(net707)
);

sky130_fd_sc_hd__xor2_2 merge844(
.A(net653),
.B(net632),
.X(net708)
);

sky130_fd_sc_hd__xnor2_2 merge845(
.A(net585),
.B(net573),
.Y(net709)
);

sky130_fd_sc_hd__xor2_1 merge846(
.A(net127),
.B(net658),
.X(net710)
);

sky130_fd_sc_hd__xnor2_4 merge847(
.A(net665),
.B(net679),
.Y(net711)
);

sky130_fd_sc_hd__xnor2_4 merge848(
.A(net255),
.B(net261),
.Y(net712)
);

sky130_fd_sc_hd__xor2_4 merge849(
.A(net283),
.B(net285),
.X(net713)
);

sky130_fd_sc_hd__xnor2_1 merge850(
.A(net310),
.B(net318),
.Y(net714)
);

sky130_fd_sc_hd__xnor2_4 merge851(
.A(net430),
.B(net304),
.Y(net715)
);

sky130_fd_sc_hd__xor2_4 merge852(
.A(net238),
.B(net668),
.X(net716)
);

sky130_fd_sc_hd__xnor2_4 merge853(
.A(net262),
.B(net663),
.Y(net717)
);

sky130_fd_sc_hd__dfrtp_2 merge854(
.D(net709),
.RESET_B(net685),
.CLK(clk),
.Q(net718)
);

sky130_fd_sc_hd__dfrtp_4 merge855(
.D(net674),
.RESET_B(net176),
.CLK(clk),
.Q(net719)
);

sky130_fd_sc_hd__xor2_1 merge856(
.A(net433),
.B(net532),
.X(net720)
);

sky130_fd_sc_hd__dfsbp_1 merge857(
.D(net151),
.SET_B(net710),
.CLK(clk),
.Q(net722),
.Q_N(net721)
);

sky130_fd_sc_hd__xnor2_4 merge858(
.A(net324),
.B(net323),
.Y(net723)
);

sky130_fd_sc_hd__xor2_1 merge859(
.A(net535),
.B(net321),
.X(net724)
);

sky130_fd_sc_hd__xnor2_1 merge860(
.A(net636),
.B(net640),
.Y(net725)
);

sky130_fd_sc_hd__xnor2_4 merge861(
.A(net631),
.B(net627),
.Y(net726)
);

sky130_fd_sc_hd__xor2_2 merge862(
.A(net639),
.B(net708),
.X(net727)
);

sky130_fd_sc_hd__xor2_1 merge863(
.A(net656),
.B(net678),
.X(net728)
);

sky130_fd_sc_hd__dfsbp_2 merge864(
.D(net723),
.SET_B(net713),
.CLK(clk),
.Q(out13),
.Q_N(net729)
);

sky130_fd_sc_hd__xor2_1 merge865(
.A(net492),
.B(net619),
.X(net730)
);

sky130_fd_sc_hd__dfstp_1 merge866(
.D(net730),
.SET_B(net672),
.CLK(clk),
.Q(net731)
);

sky130_fd_sc_hd__dfstp_2 merge867(
.D(net714),
.SET_B(net692),
.CLK(clk),
.Q(out42)
);

sky130_fd_sc_hd__xor2_1 merge868(
.A(net539),
.B(net652),
.X(net732)
);

sky130_fd_sc_hd__dfstp_4 merge869(
.D(net387),
.SET_B(net609),
.CLK(clk),
.Q(net733)
);

sky130_fd_sc_hd__dlrbn_1 merge870(
.D(net495),
.RESET_B(net702),
.GATE_N(clk),
.Q(net735),
.Q_N(net734)
);

sky130_fd_sc_hd__dlrbn_2 merge871(
.D(net696),
.RESET_B(net148),
.GATE_N(clk),
.Q(net737),
.Q_N(net736)
);

sky130_fd_sc_hd__xnor2_4 merge872(
.A(net654),
.B(net319),
.Y(net738)
);

sky130_fd_sc_hd__dlrbp_1 merge873(
.D(net669),
.RESET_B(net676),
.GATE(clk),
.Q(net740),
.Q_N(net739)
);

sky130_fd_sc_hd__dlrbp_2 merge874(
.D(net684),
.RESET_B(net701),
.GATE(clk),
.Q(net742),
.Q_N(net741)
);

sky130_fd_sc_hd__dlrtn_1 merge875(
.D(net671),
.RESET_B(net664),
.GATE_N(clk),
.Q(net743)
);

sky130_fd_sc_hd__dlrtn_2 merge876(
.D(net715),
.RESET_B(net682),
.GATE_N(clk),
.Q(net744)
);

sky130_fd_sc_hd__dlrtn_4 merge877(
.D(net681),
.RESET_B(net673),
.GATE_N(clk),
.Q(net745)
);

sky130_fd_sc_hd__dlrtp_1 merge878(
.D(net657),
.RESET_B(net466),
.GATE(clk),
.Q(net746)
);

sky130_fd_sc_hd__dlrtp_2 merge879(
.D(net686),
.RESET_B(net688),
.GATE(clk),
.Q(net747)
);

sky130_fd_sc_hd__dlrtp_4 merge880(
.Q(net388),
.RESET_B(net706),
.GATE(clk)
);

sky130_fd_sc_hd__edfxbp_1 merge881(
.D(net726),
.DE(net660),
.CLK(clk),
.Q(out11),
.Q_N(net749)
);

sky130_fd_sc_hd__xnor2_1 merge882(
.A(net634),
.B(net651),
.Y(net750)
);

sky130_fd_sc_hd__edfxtp_1 merge883(
.D(net195),
.DE(net154),
.CLK(clk),
.Q(net751)
);

sky130_fd_sc_hd__sdlclkp_1 merge884(
.GATE(net476),
.SCE(net724),
.CLK(clk),
.GCLK(out22)
);

sky130_fd_sc_hd__xor2_1 merge885(
.A(net601),
.B(net473),
.X(net752)
);

sky130_fd_sc_hd__xnor2_2 merge886(
.A(net317),
.B(net313),
.Y(net753)
);

sky130_fd_sc_hd__sdlclkp_2 merge887(
.GATE(net720),
.SCE(net662),
.CLK(clk),
.GCLK(out35)
);

sky130_fd_sc_hd__xnor2_1 merge888(
.A(net638),
.B(net635),
.Y(net754)
);

sky130_fd_sc_hd__sdlclkp_4 merge889(
.GATE(net252),
.SCE(net705),
.CLK(clk),
.GCLK(net755)
);

sky130_fd_sc_hd__dfrbp_1 merge890(
.D(net280),
.RESET_B(net400),
.CLK(clk),
.Q(net757),
.Q_N(net756)
);

sky130_fd_sc_hd__xnor2_2 merge891(
.A(net650),
.B(net637),
.Y(net758)
);

sky130_fd_sc_hd__xor2_4 merge892(
.A(net647),
.B(net646),
.X(net759)
);

sky130_fd_sc_hd__dfrbp_2 merge893(
.D(net642),
.RESET_B(net527),
.CLK(clk),
.Q(net761),
.Q_N(net760)
);

sky130_fd_sc_hd__dfrtn_1 merge894(
.D(net704),
.RESET_B(net732),
.CLK_N(clk),
.Q(out30)
);

sky130_fd_sc_hd__dfrtp_1 merge895(
.D(net597),
.RESET_B(net759),
.CLK(clk),
.Q(out19)
);

sky130_fd_sc_hd__dfrtp_2 merge896(
.D(net689),
.RESET_B(net758),
.CLK(clk),
.Q(out5)
);

sky130_fd_sc_hd__xor2_2 merge897(
.A(net541),
.B(net531),
.X(net762)
);

sky130_fd_sc_hd__dfrtp_4 merge898(
.D(net690),
.RESET_B(net282),
.CLK(clk),
.Q(out44)
);

sky130_fd_sc_hd__dfsbp_1 merge899(
.D(net284),
.SET_B(net753),
.CLK(clk),
.Q(out53),
.Q_N(net763)
);

sky130_fd_sc_hd__dfsbp_2 merge900(
.D(net305),
.SET_B(net728),
.CLK(clk),
.Q(net765),
.Q_N(net764)
);

sky130_fd_sc_hd__dfstp_1 merge901(
.D(net659),
.SET_B(net628),
.CLK(clk),
.Q(net766)
);

sky130_fd_sc_hd__dfstp_2 merge902(
.D(net691),
.SET_B(net707),
.CLK(clk),
.Q(net767)
);

sky130_fd_sc_hd__dfstp_4 merge903(
.D(net499),
.SET_B(net700),
.CLK(clk),
.Q(net768)
);

sky130_fd_sc_hd__dlrbn_1 merge904(
.D(net582),
.RESET_B(net754),
.GATE_N(clk),
.Q(net770),
.Q_N(net769)
);

sky130_fd_sc_hd__dlrbn_2 merge905(
.D(net677),
.RESET_B(net441),
.GATE_N(clk),
.Q(net772),
.Q_N(net771)
);

sky130_fd_sc_hd__dlrbp_1 merge906(
.D(net221),
.RESET_B(net306),
.GATE(clk),
.Q(net774),
.Q_N(net773)
);

sky130_fd_sc_hd__dlrbp_2 merge907(
.D(net750),
.RESET_B(net727),
.GATE(clk),
.Q(out1),
.Q_N(net775)
);

sky130_fd_sc_hd__dlrtn_1 merge908(
.D(net725),
.RESET_B(net626),
.GATE_N(clk),
.Q(net776)
);

sky130_fd_sc_hd__dlrtn_2 merge909(
.D(net693),
.RESET_B(net453),
.GATE_N(clk),
.Q(net777)
);

sky130_fd_sc_hd__dlrtn_4 merge910(
.D(net474),
.RESET_B(net416),
.GATE_N(clk),
.Q(net778)
);

sky130_fd_sc_hd__dlrtp_1 merge911(
.D(net611),
.RESET_B(net687),
.GATE(clk),
.Q(net779)
);

sky130_fd_sc_hd__dlrtp_2 merge912(
.D(net698),
.RESET_B(net610),
.GATE(clk),
.Q(net780)
);

sky130_fd_sc_hd__dlrtp_4 merge913(
.D(net242),
.RESET_B(net716),
.GATE(clk),
.Q(net781)
);

sky130_fd_sc_hd__edfxbp_1 merge914(
.D(net506),
.DE(net762),
.CLK(clk),
.Q(net782),
.Q_N(out17)
);

sky130_fd_sc_hd__edfxtp_1 merge915(
.D(net712),
.DE(net717),
.CLK(clk),
.Q(net783)
);

sky130_fd_sc_hd__sdlclkp_1 merge916(
.GATE(net699),
.SCE(net516),
.CLK(clk),
.GCLK(out21)
);

sky130_fd_sc_hd__sdlclkp_2 merge917(
.GATE(net560),
.SCE(net584),
.CLK(clk),
.GCLK(net784)
);

sky130_fd_sc_hd__sdlclkp_4 merge918(
.GATE(net620),
.SCE(net623),
.CLK(clk),
.GCLK(net785)
);

sky130_fd_sc_hd__dfrbp_1 merge919(
.D(net576),
.RESET_B(net752),
.CLK(clk),
.Q(net787),
.Q_N(net786)
);

sky130_fd_sc_hd__dfrbp_2 merge920(
.D(net711),
.RESET_B(net738),
.CLK(clk),
.Q(net788),
.Q_N(out20)
);

sky130_fd_sc_hd__dfxbp_1 s921(
.D(net58),
.CLK(clk),
.Q(net790),
.Q_N(net789)
);

sky130_fd_sc_hd__dfxbp_2 s922(
.D(net63),
.CLK(clk),
.Q(net792),
.Q_N(net791)
);

sky130_fd_sc_hd__dfxtp_1 s923(
.D(net64),
.CLK(clk),
.Q(net793)
);

sky130_fd_sc_hd__dfxtp_2 s924(
.D(net66),
.CLK(clk),
.Q(out34)
);

sky130_fd_sc_hd__dfxtp_4 s925(
.D(net133),
.CLK(clk),
.Q(net794)
);

sky130_fd_sc_hd__dlclkp_1 s926(
.GATE(net168),
.CLK(clk),
.GCLK(out2)
);

sky130_fd_sc_hd__dlclkp_2 s927(
.GATE(net189),
.CLK(clk),
.GCLK(net795)
);

sky130_fd_sc_hd__dlclkp_4 s928(
.GATE(net196),
.CLK(clk),
.GCLK(net796)
);

sky130_fd_sc_hd__dlxbn_1 s929(
.D(net215),
.GATE_N(clk),
.Q(net798),
.Q_N(net797)
);

sky130_fd_sc_hd__dlxbn_2 s930(
.D(net260),
.GATE_N(clk),
.Q(net800),
.Q_N(net799)
);

sky130_fd_sc_hd__dlxbp_1 s931(
.D(net338),
.GATE(clk),
.Q(net802),
.Q_N(net801)
);

sky130_fd_sc_hd__dlxtn_1 s932(
.D(net376),
.GATE_N(clk),
.Q(net803)
);

sky130_fd_sc_hd__dlxtn_2 s933(
.D(net382),
.GATE_N(clk),
.Q(net804)
);

sky130_fd_sc_hd__dlxtn_4 s934(
.D(net383),
.GATE_N(clk),
.Q(net805)
);

sky130_fd_sc_hd__dlxtp_1 s935(
.D(net389),
.GATE(clk),
.Q(net806)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s936(
.D(net398),
.SLEEP_B(clk),
.Q(net807)
);

sky130_fd_sc_hd__dfxbp_1 s937(
.D(net427),
.CLK(clk),
.Q(net809),
.Q_N(net808)
);

sky130_fd_sc_hd__dfxbp_2 s938(
.D(net520),
.CLK(clk),
.Q(out9),
.Q_N(net810)
);

sky130_fd_sc_hd__dfxtp_1 s939(
.D(net523),
.CLK(clk),
.Q(net811)
);

sky130_fd_sc_hd__dfxtp_2 s940(
.D(net537),
.CLK(clk),
.Q(net812)
);

sky130_fd_sc_hd__dfxtp_4 s941(
.D(net563),
.CLK(clk),
.Q(net813)
);

sky130_fd_sc_hd__dlclkp_1 s942(
.GATE(net586),
.CLK(clk),
.GCLK(net814)
);

sky130_fd_sc_hd__dlclkp_2 s943(
.GATE(net589),
.CLK(clk),
.GCLK(net815)
);

sky130_fd_sc_hd__dlclkp_4 s944(
.GATE(net598),
.CLK(clk),
.GCLK(net816)
);

sky130_fd_sc_hd__dlxbn_1 s945(
.D(net605),
.GATE_N(clk),
.Q(net818),
.Q_N(net817)
);

sky130_fd_sc_hd__dlxbn_2 s946(
.D(net606),
.GATE_N(clk),
.Q(net820),
.Q_N(net819)
);

sky130_fd_sc_hd__dlxbp_1 s947(
.D(net607),
.GATE(clk),
.Q(net822),
.Q_N(net821)
);

sky130_fd_sc_hd__dlxtn_1 s948(
.D(net608),
.GATE_N(clk),
.Q(net823)
);

sky130_fd_sc_hd__dlxtn_2 s949(
.D(net618),
.GATE_N(clk),
.Q(net824)
);

sky130_fd_sc_hd__dlxtn_4 s950(
.D(net645),
.GATE_N(clk),
.Q(net825)
);

sky130_fd_sc_hd__dlxtp_1 s951(
.D(net648),
.GATE(clk),
.Q(out3)
);


endmodule
