module netlist_1 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input in52,
	input in53,
	input in54,
	input in55,
	input in56,
	input in57,
	input in58,
	input in59,
	input in60,
	input in61,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51,
	output out52,
	output out53,
	output out54,
	output out55,
	output out56,
	output out57,
	output out58,
	output out59,
	output out60,
	output out61
);


wire clk;
wire net893;
wire net892;
wire net890;
wire net889;
wire net885;
wire net882;
wire net881;
wire net880;
wire net878;
wire net877;
wire net887;
wire net875;
wire net871;
wire out20;
wire net866;
wire net865;
wire net864;
wire net863;
wire net862;
wire net860;
wire net857;
wire net854;
wire net853;
wire net851;
wire net850;
wire net849;
wire net848;
wire net846;
wire net844;
wire net842;
wire net841;
wire net837;
wire net834;
wire net833;
wire net832;
wire net831;
wire net829;
wire net827;
wire net825;
wire net843;
wire net823;
wire net822;
wire net821;
wire net820;
wire net819;
wire out43;
wire net818;
wire net817;
wire net816;
wire net815;
wire net814;
wire net813;
wire net812;
wire net811;
wire net810;
wire net807;
wire out2;
wire net805;
wire net804;
wire net802;
wire net801;
wire net800;
wire net795;
wire out37;
wire net793;
wire net792;
wire net791;
wire out40;
wire net789;
wire out24;
wire net787;
wire net786;
wire net785;
wire net784;
wire net808;
wire net781;
wire net780;
wire net777;
wire net869;
wire net776;
wire net775;
wire net774;
wire net773;
wire net772;
wire net771;
wire net770;
wire net769;
wire out35;
wire net766;
wire net765;
wire net764;
wire net763;
wire net762;
wire net759;
wire net755;
wire net754;
wire net753;
wire net752;
wire net751;
wire net750;
wire net748;
wire net790;
wire net747;
wire net745;
wire out45;
wire net744;
wire net743;
wire net741;
wire net740;
wire net739;
wire net738;
wire net735;
wire net732;
wire net731;
wire net730;
wire net729;
wire net728;
wire net726;
wire net725;
wire net724;
wire net722;
wire net720;
wire net719;
wire net717;
wire net716;
wire net715;
wire net714;
wire net712;
wire net711;
wire net708;
wire net706;
wire net705;
wire net704;
wire net703;
wire net701;
wire net699;
wire net779;
wire net698;
wire net697;
wire net696;
wire net695;
wire net694;
wire net693;
wire net692;
wire net690;
wire net895;
wire net299;
wire net688;
wire net686;
wire net684;
wire net683;
wire net503;
wire net679;
wire net671;
wire net669;
wire net668;
wire net370;
wire net667;
wire net664;
wire net659;
wire in6;
wire net656;
wire net652;
wire net622;
wire net651;
wire net304;
wire net645;
wire net641;
wire net637;
wire net632;
wire net665;
wire net631;
wire net629;
wire net74;
wire net628;
wire net3;
wire net627;
wire net447;
wire net626;
wire net624;
wire net506;
wire net623;
wire net620;
wire in49;
wire net619;
wire net879;
wire net798;
wire net46;
wire net615;
wire net100;
wire net347;
wire net288;
wire net614;
wire net165;
wire net613;
wire net20;
wire net612;
wire net638;
wire net428;
wire net610;
wire out25;
wire net608;
wire net1;
wire net424;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire net782;
wire net601;
wire net596;
wire net592;
wire net588;
wire net587;
wire in4;
wire net583;
wire net707;
wire net582;
wire net158;
wire net584;
wire net581;
wire net336;
wire net579;
wire net577;
wire net576;
wire net570;
wire net209;
wire net569;
wire in41;
wire net567;
wire net794;
wire in30;
wire net566;
wire net565;
wire net39;
wire net562;
wire net559;
wire net556;
wire net876;
wire net647;
wire net555;
wire net159;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire in55;
wire net550;
wire net867;
wire net710;
wire net544;
wire net539;
wire net534;
wire net532;
wire net271;
wire net530;
wire net617;
wire net306;
wire net537;
wire net369;
wire net528;
wire net525;
wire net523;
wire net872;
wire net520;
wire net519;
wire net516;
wire net672;
wire net514;
wire out18;
wire net78;
wire net508;
wire net721;
wire net504;
wire net224;
wire net573;
wire net499;
wire net674;
wire net496;
wire net495;
wire net494;
wire net888;
wire net179;
wire in39;
wire net453;
wire net493;
wire net788;
wire net472;
wire net492;
wire net897;
wire net479;
wire net491;
wire net295;
wire net490;
wire net489;
wire net856;
wire net487;
wire net486;
wire net478;
wire net474;
wire net473;
wire net468;
wire net540;
wire net202;
wire net465;
wire out7;
wire net462;
wire net469;
wire net471;
wire net461;
wire net546;
wire net749;
wire net460;
wire net454;
wire net44;
wire net117;
wire net689;
wire net859;
wire net858;
wire net648;
wire net452;
wire net449;
wire net448;
wire net498;
wire net700;
wire net446;
wire net680;
wire net691;
wire net88;
wire net444;
wire in59;
wire net110;
wire net442;
wire net609;
wire net440;
wire net128;
wire net439;
wire out21;
wire net147;
wire net438;
wire net797;
wire net433;
wire net432;
wire out41;
wire net419;
wire net431;
wire net430;
wire net618;
wire net429;
wire net427;
wire net809;
wire net426;
wire net673;
wire net425;
wire net423;
wire net183;
wire net531;
wire net421;
wire net52;
wire net170;
wire net420;
wire net450;
wire net418;
wire net416;
wire net415;
wire net414;
wire net276;
wire net413;
wire net330;
wire net252;
wire net412;
wire net411;
wire net826;
wire net517;
wire net677;
wire net410;
wire net409;
wire out17;
wire net685;
wire net407;
wire out19;
wire net406;
wire net662;
wire net405;
wire net836;
wire net607;
wire net526;
wire net404;
wire net29;
wire net403;
wire net383;
wire net663;
wire net402;
wire net106;
wire net572;
wire net401;
wire net847;
wire net399;
wire net398;
wire net476;
wire net855;
wire net396;
wire out3;
wire net172;
wire net395;
wire net391;
wire net884;
wire net443;
wire net557;
wire net345;
wire net527;
wire net488;
wire net390;
wire out5;
wire net646;
wire net389;
wire net513;
wire out14;
wire net501;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net184;
wire net131;
wire net380;
wire net379;
wire net260;
wire net616;
wire net378;
wire net543;
wire net38;
wire net377;
wire net376;
wire net625;
wire net373;
wire net598;
wire net374;
wire net676;
wire net861;
wire net372;
wire net371;
wire net368;
wire net367;
wire net366;
wire net365;
wire net364;
wire net363;
wire net360;
wire net397;
wire net357;
wire net356;
wire net510;
wire net355;
wire out13;
wire net590;
wire net507;
wire net351;
wire net746;
wire net350;
wire net547;
wire net511;
wire net451;
wire net13;
wire net343;
wire net89;
wire net666;
wire net340;
wire net339;
wire net337;
wire net458;
wire net538;
wire net244;
wire net334;
wire net333;
wire net332;
wire net331;
wire net328;
wire net327;
wire net119;
wire net325;
wire net324;
wire net321;
wire net535;
wire net320;
wire net542;
wire net139;
wire net318;
wire out31;
wire net316;
wire out9;
wire net335;
wire net315;
wire net313;
wire net505;
wire net199;
wire out27;
wire net294;
wire net319;
wire net312;
wire net309;
wire net742;
wire net308;
wire net352;
wire net845;
wire net307;
wire net305;
wire net291;
wire net303;
wire net301;
wire net298;
wire net296;
wire in24;
wire net358;
wire net127;
wire net293;
wire net594;
wire out39;
wire net292;
wire net500;
wire net445;
wire net230;
wire out22;
wire net201;
wire net422;
wire net289;
wire net595;
wire net384;
wire net482;
wire in25;
wire net589;
wire net278;
wire net761;
wire net274;
wire net643;
wire net273;
wire net272;
wire net114;
wire net270;
wire in17;
wire net267;
wire net644;
wire net266;
wire net459;
wire net463;
wire net0;
wire net297;
wire net408;
wire net475;
wire net280;
wire net102;
wire net799;
wire net151;
wire net275;
wire net264;
wire net657;
wire net591;
wire net196;
wire net262;
wire net217;
wire net261;
wire net21;
wire net257;
wire net62;
wire net109;
wire net254;
wire net203;
wire net253;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire net660;
wire net838;
wire net359;
wire out28;
wire net417;
wire net302;
wire out8;
wire in26;
wire net661;
wire net194;
wire net241;
wire in29;
wire net240;
wire out42;
wire net238;
wire out10;
wire net142;
wire net234;
wire net232;
wire out12;
wire net226;
wire out32;
wire net568;
wire net375;
wire net223;
wire net524;
wire net575;
wire net382;
wire net852;
wire net548;
wire net259;
wire net222;
wire net31;
wire net219;
wire net578;
wire net210;
wire net326;
wire net213;
wire net208;
wire out16;
wire net188;
wire net891;
wire net207;
wire net649;
wire net205;
wire net678;
wire net633;
wire net122;
wire net197;
wire net840;
wire net483;
wire net193;
wire net192;
wire net737;
wire net190;
wire net630;
wire in20;
wire net874;
wire net189;
wire net246;
wire net783;
wire net186;
wire net152;
wire net126;
wire net113;
wire net284;
wire net655;
wire net563;
wire net464;
wire net549;
wire net182;
wire net310;
wire net180;
wire in8;
wire net30;
wire out36;
wire net342;
wire net17;
wire net886;
wire net437;
wire out44;
wire out58;
wire net580;
wire net133;
wire net175;
wire out56;
wire out38;
wire net80;
wire net173;
wire net521;
wire net353;
wire in37;
wire net518;
wire net381;
wire net218;
wire net300;
wire net169;
wire net828;
wire net485;
wire net344;
wire net168;
wire net153;
wire net286;
wire net167;
wire net509;
wire net58;
wire net221;
wire net166;
wire net269;
wire net97;
wire net434;
wire net204;
wire net200;
wire net621;
wire net162;
wire out60;
wire net497;
wire net161;
wire net285;
wire net160;
wire net636;
wire net311;
wire net441;
wire out15;
wire net150;
wire net149;
wire net148;
wire net178;
wire net239;
wire net144;
wire net322;
wire net758;
wire net143;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net806;
wire net561;
wire out29;
wire net137;
wire net136;
wire net456;
wire net868;
wire net135;
wire net255;
wire net157;
wire net177;
wire net349;
wire out51;
wire out48;
wire net134;
wire net250;
wire net225;
wire net132;
wire net130;
wire net242;
wire net124;
wire net642;
wire net268;
wire in7;
wire net756;
wire net400;
wire net82;
wire net870;
wire net2;
wire net123;
wire net481;
wire net120;
wire net392;
wire net164;
wire net687;
wire net282;
wire net71;
wire net229;
wire in43;
wire net108;
wire net107;
wire out33;
wire net41;
wire net8;
wire net104;
wire in12;
wire net894;
wire net103;
wire out26;
wire net99;
wire net348;
wire net341;
wire in52;
wire net6;
wire net457;
wire out50;
wire net96;
wire net466;
wire net118;
wire net94;
wire net90;
wire net803;
wire net174;
wire net277;
wire net639;
wire net81;
wire in10;
wire net156;
wire net361;
wire net115;
wire net670;
wire in18;
wire net27;
wire net34;
wire net585;
wire net79;
wire out6;
wire net231;
wire net329;
wire net212;
wire net653;
wire in5;
wire net14;
wire net77;
wire net600;
wire net236;
wire net76;
wire in42;
wire net354;
wire in38;
wire net736;
wire net198;
wire net467;
wire net101;
wire net9;
wire net75;
wire net42;
wire net91;
wire out4;
wire net873;
wire net571;
wire net73;
wire net60;
wire net564;
wire net154;
wire net84;
wire net237;
wire net682;
wire in46;
wire net85;
wire net72;
wire net116;
wire net69;
wire net67;
wire in31;
wire net129;
wire net65;
wire net98;
wire net522;
wire net436;
wire net541;
wire net323;
wire net15;
wire net279;
wire net64;
wire net63;
wire net681;
wire net61;
wire net512;
wire net18;
wire out34;
wire net59;
wire net248;
wire net477;
wire net228;
wire net675;
wire net56;
wire net55;
wire net214;
wire net53;
wire in48;
wire net640;
wire net50;
wire out49;
wire out61;
wire net597;
wire net185;
wire net155;
wire net338;
wire net599;
wire net112;
wire net195;
wire out52;
wire net650;
wire net560;
wire net45;
wire net502;
wire net235;
wire net830;
wire net49;
wire in50;
wire net215;
wire net484;
wire net346;
wire net4;
wire net43;
wire net187;
wire in13;
wire net586;
wire net533;
wire net796;
wire net32;
wire net125;
wire net19;
wire in15;
wire net896;
wire net727;
wire net163;
wire in19;
wire net702;
wire net70;
wire net48;
wire net28;
wire net92;
wire net713;
wire net25;
wire out59;
wire in0;
wire net709;
wire net24;
wire out47;
wire net290;
wire net227;
wire net258;
wire net176;
wire net839;
wire out23;
wire net470;
wire in33;
wire net33;
wire net824;
wire net233;
wire net40;
wire in60;
wire net435;
wire net760;
wire net23;
wire net26;
wire net16;
wire net558;
wire in1;
wire net265;
wire net778;
wire net22;
wire net263;
wire net5;
wire net206;
wire in58;
wire in61;
wire net757;
wire in56;
wire net733;
wire net171;
wire in23;
wire in57;
wire net281;
wire net54;
wire in54;
wire in53;
wire net835;
wire out11;
wire net138;
wire net145;
wire net211;
wire in35;
wire in34;
wire net593;
wire in45;
wire net393;
wire net256;
wire net87;
wire net181;
wire net7;
wire out1;
wire out54;
wire net574;
wire net216;
wire net455;
wire in28;
wire in44;
wire net883;
wire in32;
wire net47;
wire net12;
wire in27;
wire in9;
wire net654;
wire net723;
wire net611;
wire net515;
wire net362;
wire in16;
wire net191;
wire out46;
wire net35;
wire net220;
wire in22;
wire net68;
wire in14;
wire net529;
wire in21;
wire net57;
wire net480;
wire net86;
wire net317;
wire in51;
wire net93;
wire in47;
wire in2;
wire net718;
wire net658;
wire net105;
wire in11;
wire net51;
wire out30;
wire in36;
wire net767;
wire net111;
wire net536;
wire net37;
wire net36;
wire net95;
wire net121;
wire net146;
wire net734;
wire net251;
wire net768;
wire net11;
wire net394;
wire net314;
wire in3;
sky130_fd_sc_hd__mux4_2 c62(
.A0(in46),
.A1(in56),
.A2(in51),
.A3(in23),
.S0(in52),
.S1(net3),
.X(net0)
);

sky130_fd_sc_hd__mux4_4 c63(
.A0(in60),
.A1(in49),
.A2(in58),
.A3(in24),
.S0(in47),
.S1(in56),
.X(net1)
);

sky130_fd_sc_hd__mux4_1 c64(
.A0(in55),
.A1(in59),
.A2(in52),
.A3(net1),
.S0(in46),
.S1(net3),
.X(net2)
);

sky130_fd_sc_hd__a2111oi_1 c65(
.A1(in24),
.A2(in36),
.B1(in23),
.C1(in20),
.D1(in29),
.Y(net3)
);

sky130_fd_sc_hd__nand2_4 c66(
.A(in54),
.B(in56),
.Y(net4)
);

sky130_fd_sc_hd__nor2_2 c67(
.A(in48),
.B(in29),
.Y(net5)
);

sky130_fd_sc_hd__nor2b_4 c68(
.A(in58),
.B_N(in57),
.Y(net6)
);

sky130_fd_sc_hd__and2_4 c69(
.A(net6),
.B(in27),
.X(net7)
);

sky130_fd_sc_hd__o2111a_1 c70(
.A1(in46),
.A2(net0),
.B1(in51),
.C1(in36),
.D1(net5),
.X(net8)
);

sky130_fd_sc_hd__and3b_2 c71(
.A_N(in56),
.B(in49),
.C(in47),
.X(net9)
);

sky130_fd_sc_hd__nand2_4 c72(
.A(net7),
.B(in58),
.Y(net10)
);

sky130_fd_sc_hd__nor3b_4 c73(
.A(in44),
.B(in53),
.C_N(net2),
.Y(net11)
);

sky130_fd_sc_hd__and2b_2 c74(
.A_N(in49),
.B(net7),
.X(net12)
);

sky130_fd_sc_hd__nand3_2 c75(
.A(net9),
.B(net4),
.C(net5),
.Y(net13)
);

sky130_fd_sc_hd__and2_1 c76(
.A(net6),
.B(net13),
.X(net14)
);

sky130_fd_sc_hd__mux4_2 c77(
.A0(in51),
.A1(net10),
.A2(net12),
.A3(in7),
.S0(net7),
.S1(net14),
.X(net15)
);

sky130_fd_sc_hd__clkbuf_4 c78(
.A(net644),
.X(net16)
);

sky130_fd_sc_hd__or2b_4 c79(
.A(in53),
.B_N(in25),
.X(net17)
);

sky130_fd_sc_hd__or4bb_2 c80(
.A(net4),
.B(net17),
.C_N(net16),
.D_N(net710),
.X(net18)
);

sky130_fd_sc_hd__buf_6 c81(
.A(net644),
.X(net19)
);

sky130_fd_sc_hd__clkbuf_8 c82(
.A(net710),
.X(net20)
);

sky130_fd_sc_hd__sdfrbp_1 c83(
.D(net11),
.RESET_B(net20),
.SCD(net16),
.SCE(net710),
.CLK(clk),
.Q(net22),
.Q_N(net21)
);

sky130_fd_sc_hd__clkinv_1 c84(
.A(net746),
.Y(net23)
);

sky130_fd_sc_hd__mux4_1 c85(
.A0(net11),
.A1(net14),
.A2(net23),
.A3(net17),
.S0(net22),
.S1(net5),
.X(net24)
);

sky130_fd_sc_hd__or4bb_4 c86(
.A(net17),
.B(net16),
.C_N(net23),
.D_N(net4),
.X(net25)
);

sky130_fd_sc_hd__mux4_2 c87(
.A0(net20),
.A1(in51),
.A2(net25),
.A3(net23),
.S0(net11),
.S1(net17),
.X(net26)
);

sky130_fd_sc_hd__inv_1 c88(
.A(net718),
.Y(net27)
);

sky130_fd_sc_hd__nand2b_2 c89(
.A_N(net0),
.B(net9),
.Y(net28)
);

sky130_fd_sc_hd__buf_12 c90(
.A(net744),
.X(net29)
);

sky130_fd_sc_hd__or3_4 c91(
.A(net0),
.B(net27),
.C(net821),
.X(net30)
);

sky130_fd_sc_hd__or3_4 c92(
.A(net9),
.B(in54),
.C(net823),
.X(net31)
);

sky130_fd_sc_hd__clkbuf_8 c93(
.A(net718),
.X(net32)
);

sky130_fd_sc_hd__and2b_1 c94(
.A_N(in29),
.B(net821),
.X(net33)
);

sky130_fd_sc_hd__dlygate4sd1_1 c95(
.A(net744),
.X(out49)
);

sky130_fd_sc_hd__and2_2 c96(
.A(out49),
.B(net823),
.X(net34)
);

sky130_fd_sc_hd__or3_1 c97(
.A(net29),
.B(in57),
.C(net820),
.X(net35)
);

sky130_fd_sc_hd__and3_2 c98(
.A(net31),
.B(in61),
.C(net33),
.X(net36)
);

sky130_fd_sc_hd__clkinv_8 c99(
.A(net779),
.Y(net37)
);

sky130_fd_sc_hd__and3b_2 c100(
.A_N(net34),
.B(net37),
.C(net7),
.X(net38)
);

sky130_fd_sc_hd__buf_16 c101(
.A(net779),
.X(net39)
);

sky130_fd_sc_hd__or3_4 c102(
.A(net33),
.B(net37),
.C(net29),
.X(net40)
);

sky130_fd_sc_hd__or4bb_4 c103(
.A(net36),
.B(net35),
.C_N(net40),
.D_N(net37),
.X(net41)
);

sky130_fd_sc_hd__sdfbbn_1 c104(
.D(in36),
.RESET_B(net19),
.SCD(net36),
.SCE(net38),
.SET_B(net718),
.CLK_N(clk),
.Q(out23),
.Q_N(net42)
);

sky130_fd_sc_hd__mux4_1 c105(
.A0(net10),
.A1(net32),
.A2(net29),
.A3(net35),
.S0(net36),
.S1(net822),
.X(net43)
);

sky130_fd_sc_hd__or4bb_2 c106(
.A(net22),
.B(out49),
.C_N(net42),
.D_N(net824),
.X(net44)
);

sky130_fd_sc_hd__mux4_1 c107(
.A0(net19),
.A1(net31),
.A2(net35),
.A3(net22),
.S0(net718),
.S1(net824),
.X(net45)
);

sky130_fd_sc_hd__sdfrbp_2 c108(
.D(net45),
.RESET_B(net35),
.SCD(out23),
.SCE(net824),
.CLK(clk),
.Q(out22),
.Q_N(net46)
);

sky130_fd_sc_hd__mux4_2 c109(
.A0(net38),
.A1(net45),
.A2(net44),
.A3(net42),
.S0(net28),
.S1(net824),
.X(net47)
);

sky130_fd_sc_hd__buf_2 c110(
.A(net656),
.X(net48)
);

sky130_fd_sc_hd__inv_4 c111(
.A(net656),
.Y(net49)
);

sky130_fd_sc_hd__nor2_4 c112(
.A(in18),
.B(in14),
.Y(out61)
);

sky130_fd_sc_hd__or2_4 c113(
.A(out61),
.B(net19),
.X(net50)
);

sky130_fd_sc_hd__or4bb_2 c114(
.A(in57),
.B(net49),
.C_N(net19),
.D_N(net28),
.X(net51)
);

sky130_fd_sc_hd__nand2_1 c115(
.A(in45),
.B(net49),
.Y(net52)
);

sky130_fd_sc_hd__and2_2 c116(
.A(net5),
.B(net49),
.X(net53)
);

sky130_fd_sc_hd__buf_12 c117(
.A(net726),
.X(net54)
);

sky130_fd_sc_hd__or2b_2 c118(
.A(net52),
.B_N(net46),
.X(net55)
);

sky130_fd_sc_hd__or2_1 c119(
.A(net19),
.B(net48),
.X(out26)
);

sky130_fd_sc_hd__a2111oi_4 c120(
.A1(net32),
.A2(in57),
.B1(net49),
.C1(net44),
.D1(out26),
.Y(out54)
);

sky130_fd_sc_hd__nor2_4 c121(
.A(net37),
.B(net19),
.Y(out29)
);

sky130_fd_sc_hd__and2_0 c122(
.A(net48),
.B(out26),
.X(net56)
);

sky130_fd_sc_hd__or4bb_1 c123(
.A(net56),
.B(net49),
.C_N(out26),
.D_N(net52),
.X(net57)
);

sky130_fd_sc_hd__or3b_2 c124(
.A(net35),
.B(out26),
.C_N(net825),
.X(net58)
);

sky130_fd_sc_hd__nand2b_4 c125(
.A_N(net44),
.B(out26),
.Y(net59)
);

sky130_fd_sc_hd__nand2_1 c126(
.A(net58),
.B(out54),
.Y(net60)
);

sky130_fd_sc_hd__buf_12 c127(
.A(net726),
.X(net61)
);

sky130_fd_sc_hd__sdfrtn_1 c128(
.D(net59),
.RESET_B(net58),
.SCD(net57),
.SCE(net49),
.CLK_N(clk),
.Q(out50)
);

sky130_fd_sc_hd__or2b_1 c129(
.A(net34),
.B_N(out50),
.X(net62)
);

sky130_fd_sc_hd__or4bb_2 c130(
.A(net53),
.B(out29),
.C_N(out50),
.D_N(out61),
.X(net63)
);

sky130_fd_sc_hd__sdfrtp_1 c131(
.D(net63),
.RESET_B(net59),
.SCD(out26),
.SCE(net19),
.CLK(clk),
.Q(out52)
);

sky130_fd_sc_hd__and3b_2 c132(
.A_N(in3),
.B(in16),
.C(in20),
.X(net64)
);

sky130_fd_sc_hd__nand2_2 c133(
.A(in5),
.B(in16),
.Y(net65)
);

sky130_fd_sc_hd__and3b_2 c134(
.A_N(in21),
.B(in18),
.C(in3),
.X(net66)
);

sky130_fd_sc_hd__and2b_4 c135(
.A_N(in19),
.B(in21),
.X(net67)
);

sky130_fd_sc_hd__nand3b_2 c136(
.A_N(in12),
.B(in17),
.C(net66),
.Y(net68)
);

sky130_fd_sc_hd__or3b_2 c137(
.A(net66),
.B(net67),
.C_N(net68),
.X(net69)
);

sky130_fd_sc_hd__and3_1 c138(
.A(net65),
.B(net68),
.C(in6),
.X(net70)
);

sky130_fd_sc_hd__and2b_4 c139(
.A_N(in13),
.B(in0),
.X(net71)
);

sky130_fd_sc_hd__mux4_2 c140(
.A0(net68),
.A1(in14),
.A2(in15),
.A3(in3),
.S0(in10),
.S1(in8),
.X(net72)
);

sky130_fd_sc_hd__and2_4 c141(
.A(in1),
.B(net71),
.X(net73)
);

sky130_fd_sc_hd__or4bb_4 c142(
.A(in0),
.B(net65),
.C_N(in20),
.D_N(in21),
.X(net74)
);

sky130_fd_sc_hd__nand3_4 c143(
.A(in6),
.B(net66),
.C(in16),
.Y(net75)
);

sky130_fd_sc_hd__clkinv_16 c144(
.A(net723),
.Y(net76)
);

sky130_fd_sc_hd__inv_16 c145(
.A(net723),
.Y(net77)
);

sky130_fd_sc_hd__mux4_1 c146(
.A0(net76),
.A1(net70),
.A2(in11),
.A3(in4),
.S0(net68),
.S1(net74),
.X(net78)
);

sky130_fd_sc_hd__or3_2 c147(
.A(net68),
.B(net74),
.C(in11),
.X(out6)
);

sky130_fd_sc_hd__a2111o_1 c148(
.A1(net77),
.A2(in0),
.B1(net75),
.C1(in17),
.D1(net72),
.X(net79)
);

sky130_fd_sc_hd__o2111ai_4 c149(
.A1(net66),
.A2(net77),
.B1(in21),
.C1(net65),
.D1(net775),
.Y(out7)
);

sky130_fd_sc_hd__mux4_2 c150(
.A0(in10),
.A1(net65),
.A2(out6),
.A3(out7),
.S0(net722),
.S1(net775),
.X(net80)
);

sky130_fd_sc_hd__mux4_2 c151(
.A0(net70),
.A1(net77),
.A2(net75),
.A3(out7),
.S0(net775),
.S1(net826),
.X(net81)
);

sky130_fd_sc_hd__mux4_1 c152(
.A0(net72),
.A1(net70),
.A2(out7),
.A3(net722),
.S0(net826),
.S1(net827),
.X(net82)
);

sky130_fd_sc_hd__mux4_4 c153(
.A0(net72),
.A1(net65),
.A2(net64),
.A3(net723),
.S0(net827),
.S1(net828),
.X(net83)
);

sky130_fd_sc_hd__nand2_2 c154(
.A(in28),
.B(in8),
.Y(net84)
);

sky130_fd_sc_hd__nand2b_1 c155(
.A_N(in8),
.B(net84),
.Y(net85)
);

sky130_fd_sc_hd__nand2_2 c156(
.A(in31),
.B(net64),
.Y(net86)
);

sky130_fd_sc_hd__or2_1 c157(
.A(in39),
.B(net85),
.X(net87)
);

sky130_fd_sc_hd__and3b_4 c158(
.A_N(in37),
.B(in34),
.C(net827),
.X(net88)
);

sky130_fd_sc_hd__or3b_4 c159(
.A(in22),
.B(net86),
.C_N(net84),
.X(net89)
);

sky130_fd_sc_hd__and2b_4 c160(
.A_N(in43),
.B(net85),
.X(net90)
);

sky130_fd_sc_hd__or2_1 c161(
.A(in32),
.B(in41),
.X(net91)
);

sky130_fd_sc_hd__sdfrtp_2 c162(
.D(net89),
.RESET_B(in15),
.SCD(net90),
.SCE(out7),
.CLK(clk),
.Q(net92)
);

sky130_fd_sc_hd__or2b_2 c163(
.A(in41),
.B_N(net92),
.X(net93)
);

sky130_fd_sc_hd__nor2_1 c164(
.A(net88),
.B(net92),
.Y(net94)
);

sky130_fd_sc_hd__clkbuf_2 c165(
.A(net775),
.X(net95)
);

sky130_fd_sc_hd__or4bb_2 c166(
.A(net90),
.B(net95),
.C_N(in8),
.D_N(net92),
.X(net96)
);

sky130_fd_sc_hd__or3_1 c167(
.A(net94),
.B(in27),
.C(net84),
.X(net97)
);

sky130_fd_sc_hd__nand2b_2 c168(
.A_N(in15),
.B(in38),
.Y(net98)
);

sky130_fd_sc_hd__and3_2 c169(
.A(net95),
.B(net94),
.C(net826),
.X(out47)
);

sky130_fd_sc_hd__mux4_1 c170(
.A0(net97),
.A1(in33),
.A2(net89),
.A3(in34),
.S0(net86),
.S1(net828),
.X(net99)
);

sky130_fd_sc_hd__nand3_4 c171(
.A(net64),
.B(net98),
.C(net85),
.Y(net100)
);

sky130_fd_sc_hd__nor3b_2 c172(
.A(net92),
.B(in37),
.C_N(net830),
.Y(net101)
);

sky130_fd_sc_hd__or4bb_2 c173(
.A(net91),
.B(net101),
.C_N(net100),
.D_N(net90),
.X(net102)
);

sky130_fd_sc_hd__clkbuf_8 c174(
.A(net775),
.X(net103)
);

sky130_fd_sc_hd__clkinv_1 c175(
.A(net755),
.Y(net104)
);

sky130_fd_sc_hd__clkbuf_1 c176(
.A(out33),
.X(net105)
);

sky130_fd_sc_hd__dlygate4sd1_1 c177(
.A(net725),
.X(net106)
);

sky130_fd_sc_hd__nor2b_2 c178(
.A(net85),
.B_N(net827),
.Y(net107)
);

sky130_fd_sc_hd__nor3_1 c179(
.A(net101),
.B(in48),
.C(in25),
.Y(net108)
);

sky130_fd_sc_hd__o2111a_1 c180(
.A1(in26),
.A2(in47),
.B1(net108),
.C1(net826),
.D1(net831),
.X(net109)
);

sky130_fd_sc_hd__inv_1 c181(
.A(out33),
.Y(net110)
);

sky130_fd_sc_hd__and2_4 c182(
.A(in26),
.B(net108),
.X(net111)
);

sky130_fd_sc_hd__clkinv_2 c183(
.A(net725),
.Y(net112)
);

sky130_fd_sc_hd__inv_8 c184(
.A(net749),
.Y(net113)
);

sky130_fd_sc_hd__clkbuf_4 c185(
.A(net755),
.X(net114)
);

sky130_fd_sc_hd__nand3b_1 c186(
.A_N(net1),
.B(in26),
.C(net112),
.Y(net115)
);

sky130_fd_sc_hd__buf_1 c187(
.A(net724),
.X(net116)
);

sky130_fd_sc_hd__nor2b_4 c188(
.A(net106),
.B_N(net112),
.Y(net117)
);

sky130_fd_sc_hd__a2111o_2 c189(
.A1(in60),
.A2(in50),
.B1(in20),
.C1(net2),
.D1(in38),
.X(net118)
);

sky130_fd_sc_hd__and3b_4 c190(
.A_N(in38),
.B(net117),
.C(net826),
.X(net119)
);

sky130_fd_sc_hd__sdfbbn_2 c191(
.D(in44),
.RESET_B(net3),
.SCD(net119),
.SCE(net118),
.SET_B(net117),
.CLK_N(clk),
.Q(net121),
.Q_N(net120)
);

sky130_fd_sc_hd__buf_8 c192(
.A(net749),
.X(net122)
);

sky130_fd_sc_hd__or3b_2 c193(
.A(net116),
.B(net119),
.C_N(in47),
.X(net123)
);

sky130_fd_sc_hd__a2111oi_4 c194(
.A1(net114),
.A2(net122),
.B1(net117),
.C1(net121),
.D1(net108),
.Y(net124)
);

sky130_fd_sc_hd__mux4_2 c195(
.A0(in23),
.A1(net123),
.A2(net124),
.A3(net108),
.S0(net107),
.S1(net93),
.X(net125)
);

sky130_fd_sc_hd__clkinv_1 c196(
.A(net771),
.Y(net126)
);

sky130_fd_sc_hd__mux4_4 c197(
.A0(net126),
.A1(net123),
.A2(net75),
.A3(net124),
.S0(net109),
.S1(net111),
.X(net127)
);

sky130_fd_sc_hd__clkinv_2 c198(
.A(net751),
.Y(net128)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c199(
.A(net751),
.X(net129)
);

sky130_fd_sc_hd__and2_4 c200(
.A(net75),
.B(net18),
.X(net130)
);

sky130_fd_sc_hd__dlygate4sd3_1 c201(
.A(net814),
.X(net131)
);

sky130_fd_sc_hd__nand2_1 c202(
.A(net20),
.B(in11),
.Y(net132)
);

sky130_fd_sc_hd__or2_1 c203(
.A(net116),
.B(net132),
.X(net133)
);

sky130_fd_sc_hd__nand2_4 c204(
.A(in27),
.B(net5),
.Y(net134)
);

sky130_fd_sc_hd__buf_2 c205(
.A(net790),
.X(net135)
);

sky130_fd_sc_hd__nand3_1 c206(
.A(net128),
.B(net75),
.C(net134),
.Y(net136)
);

sky130_fd_sc_hd__inv_16 c207(
.A(net762),
.Y(net137)
);

sky130_fd_sc_hd__inv_1 c208(
.A(net755),
.Y(net138)
);

sky130_fd_sc_hd__buf_4 c209(
.A(net762),
.X(net139)
);

sky130_fd_sc_hd__a2111o_2 c210(
.A1(net2),
.A2(net133),
.B1(net132),
.C1(net115),
.D1(net128),
.X(net140)
);

sky130_fd_sc_hd__clkinv_1 c211(
.A(net748),
.Y(net141)
);

sky130_fd_sc_hd__clkbuf_16 c212(
.A(net813),
.X(net142)
);

sky130_fd_sc_hd__sdfbbp_1 c213(
.D(net136),
.RESET_B(net128),
.SCD(net138),
.SCE(net16),
.SET_B(net131),
.CLK(clk),
.Q(net144),
.Q_N(net143)
);

sky130_fd_sc_hd__buf_2 c214(
.A(net755),
.X(net145)
);

sky130_fd_sc_hd__nand3b_2 c215(
.A_N(net141),
.B(net2),
.C(net143),
.Y(net146)
);

sky130_fd_sc_hd__o2111ai_1 c216(
.A1(net145),
.A2(net146),
.B1(net132),
.C1(net140),
.D1(net109),
.Y(net147)
);

sky130_fd_sc_hd__o2111ai_1 c217(
.A1(in7),
.A2(net145),
.B1(net131),
.C1(net142),
.D1(net143),
.Y(net148)
);

sky130_fd_sc_hd__clkbuf_4 c218(
.A(net710),
.X(net149)
);

sky130_fd_sc_hd__a2111oi_1 c219(
.A1(net149),
.A2(in7),
.B1(net130),
.C1(net148),
.D1(net832),
.Y(net150)
);

sky130_fd_sc_hd__clkinv_8 c220(
.A(net760),
.Y(net151)
);

sky130_fd_sc_hd__buf_2 c221(
.A(net760),
.X(net152)
);

sky130_fd_sc_hd__nor3_1 c222(
.A(net27),
.B(net113),
.C(net833),
.Y(net153)
);

sky130_fd_sc_hd__inv_8 c223(
.A(net762),
.Y(net154)
);

sky130_fd_sc_hd__nor3_4 c224(
.A(net139),
.B(net153),
.C(net105),
.Y(net155)
);

sky130_fd_sc_hd__or3_1 c225(
.A(net113),
.B(net106),
.C(net31),
.X(net156)
);

sky130_fd_sc_hd__sdfbbn_1 c226(
.D(net106),
.RESET_B(net39),
.SCD(net156),
.SCE(net148),
.SET_B(net824),
.CLK_N(clk),
.Q(out46),
.Q_N(net157)
);

sky130_fd_sc_hd__and3b_1 c227(
.A_N(net145),
.B(net93),
.C(net833),
.X(net158)
);

sky130_fd_sc_hd__mux4_1 c228(
.A0(net154),
.A1(net151),
.A2(net39),
.A3(net157),
.S0(net825),
.S1(net832),
.X(out15)
);

sky130_fd_sc_hd__or3b_1 c229(
.A(net154),
.B(in54),
.C_N(net158),
.X(net159)
);

sky130_fd_sc_hd__a2111oi_2 c230(
.A1(net86),
.A2(out15),
.B1(net39),
.C1(net159),
.D1(net151),
.Y(net160)
);

sky130_fd_sc_hd__sdfbbn_2 c231(
.D(net39),
.RESET_B(net158),
.SCD(net72),
.SCE(net155),
.SET_B(net148),
.CLK_N(clk),
.Q(net162),
.Q_N(net161)
);

sky130_fd_sc_hd__or4bb_1 c232(
.A(in29),
.B(net108),
.C_N(net162),
.D_N(in18),
.X(net163)
);

sky130_fd_sc_hd__a2111o_1 c233(
.A1(net40),
.A2(net155),
.B1(net162),
.C1(net39),
.D1(net157),
.X(net164)
);

sky130_fd_sc_hd__a2111o_2 c234(
.A1(net164),
.A2(net158),
.B1(net162),
.C1(net155),
.D1(net145),
.X(net165)
);

sky130_fd_sc_hd__sdfrtp_4 c235(
.D(net162),
.RESET_B(net159),
.SCD(net135),
.SCE(net734),
.CLK(clk),
.Q(out12)
);

sky130_fd_sc_hd__mux4_2 c236(
.A0(net156),
.A1(in34),
.A2(net161),
.A3(out12),
.S0(net735),
.S1(net819),
.X(net166)
);

sky130_fd_sc_hd__o2111a_2 c237(
.A1(out15),
.A2(net164),
.B1(net161),
.C1(net734),
.D1(net836),
.X(net167)
);

sky130_fd_sc_hd__mux4_2 c238(
.A0(net154),
.A1(net161),
.A2(in47),
.A3(net151),
.S0(net748),
.S1(net836),
.X(net168)
);

sky130_fd_sc_hd__a2111o_2 c239(
.A1(net168),
.A2(net164),
.B1(net161),
.C1(net748),
.D1(net824),
.X(net169)
);

sky130_fd_sc_hd__o2111ai_4 c240(
.A1(net163),
.A2(net168),
.B1(net14),
.C1(net759),
.D1(net836),
.Y(net170)
);

sky130_fd_sc_hd__mux4_1 c241(
.A0(out12),
.A1(net36),
.A2(net163),
.A3(net151),
.S0(out7),
.S1(net735),
.X(net171)
);

sky130_fd_sc_hd__buf_2 c242(
.A(out14),
.X(out25)
);

sky130_fd_sc_hd__nand2_1 c243(
.A(out46),
.B(net837),
.Y(out51)
);

sky130_fd_sc_hd__inv_4 c244(
.A(net762),
.Y(out59)
);

sky130_fd_sc_hd__and3b_4 c245(
.A_N(in14),
.B(out7),
.C(net726),
.X(net172)
);

sky130_fd_sc_hd__nand2_4 c246(
.A(net50),
.B(out12),
.Y(net173)
);

sky130_fd_sc_hd__nand3_2 c247(
.A(net49),
.B(out52),
.C(net157),
.Y(out38)
);

sky130_fd_sc_hd__and2b_4 c248(
.A_N(out50),
.B(net759),
.X(net174)
);

sky130_fd_sc_hd__a2111o_1 c249(
.A1(out52),
.A2(out26),
.B1(net825),
.C1(net836),
.D1(net837),
.X(out1)
);

sky130_fd_sc_hd__and3_4 c250(
.A(net54),
.B(net135),
.C(net829),
.X(out30)
);

sky130_fd_sc_hd__or2b_1 c251(
.A(net62),
.B_N(out26),
.X(net175)
);

sky130_fd_sc_hd__dlygate4sd3_1 c252(
.A(net748),
.X(net176)
);

sky130_fd_sc_hd__or4bb_1 c253(
.A(net159),
.B(out30),
.C_N(net176),
.D_N(net173),
.X(net177)
);

sky130_fd_sc_hd__nor2_2 c254(
.A(net135),
.B(net176),
.Y(out58)
);

sky130_fd_sc_hd__nand2b_4 c255(
.A_N(net137),
.B(net61),
.Y(net178)
);

sky130_fd_sc_hd__or2_4 c256(
.A(net174),
.B(net176),
.X(out34)
);

sky130_fd_sc_hd__nor3_1 c257(
.A(net176),
.B(out49),
.C(out61),
.Y(net179)
);

sky130_fd_sc_hd__clkbuf_1 c258(
.A(net772),
.X(out44)
);

sky130_fd_sc_hd__buf_12 c259(
.A(out14),
.X(out4)
);

sky130_fd_sc_hd__nand3_4 c260(
.A(net178),
.B(out4),
.C(net176),
.Y(out36)
);

sky130_fd_sc_hd__clkinv_16 c261(
.A(net772),
.Y(net180)
);

sky130_fd_sc_hd__mux4_4 c262(
.A0(net180),
.A1(out4),
.A2(net5),
.A3(net157),
.S0(net726),
.S1(net837),
.X(net181)
);

sky130_fd_sc_hd__mux4_4 c263(
.A0(net179),
.A1(net181),
.A2(in45),
.A3(out59),
.S0(out52),
.S1(out4),
.X(out5)
);

sky130_fd_sc_hd__clkbuf_2 c264(
.A(net728),
.X(net182)
);

sky130_fd_sc_hd__inv_2 c265(
.A(net728),
.Y(net183)
);

sky130_fd_sc_hd__nor2b_1 c266(
.A(in20),
.B_N(net71),
.Y(net184)
);

sky130_fd_sc_hd__and2b_1 c267(
.A_N(net183),
.B(in17),
.X(net185)
);

sky130_fd_sc_hd__nor2b_2 c268(
.A(net74),
.B_N(net185),
.Y(net186)
);

sky130_fd_sc_hd__clkbuf_2 c269(
.A(net728),
.X(net187)
);

sky130_fd_sc_hd__or2b_2 c270(
.A(out7),
.B_N(net184),
.X(net188)
);

sky130_fd_sc_hd__nor2_4 c271(
.A(net182),
.B(net65),
.Y(net189)
);

sky130_fd_sc_hd__clkbuf_16 c272(
.A(net780),
.X(net190)
);

sky130_fd_sc_hd__or4bb_4 c273(
.A(net188),
.B(net190),
.C_N(out7),
.D_N(net184),
.X(net191)
);

sky130_fd_sc_hd__or4bb_2 c274(
.A(net183),
.B(out7),
.C_N(net184),
.D_N(net815),
.X(net192)
);

sky130_fd_sc_hd__nand2_1 c275(
.A(net190),
.B(in14),
.Y(net193)
);

sky130_fd_sc_hd__nor3b_2 c276(
.A(net183),
.B(net189),
.C_N(net184),
.Y(net194)
);

sky130_fd_sc_hd__inv_16 c277(
.A(net768),
.Y(net195)
);

sky130_fd_sc_hd__mux4_1 c278(
.A0(net185),
.A1(net184),
.A2(net64),
.A3(net195),
.S0(out7),
.S1(net815),
.X(net196)
);

sky130_fd_sc_hd__sdfbbp_1 c279(
.D(net195),
.RESET_B(net194),
.SCD(out7),
.SCE(net189),
.SET_B(net182),
.CLK(clk),
.Q(net198),
.Q_N(net197)
);

sky130_fd_sc_hd__inv_2 c280(
.A(net768),
.Y(net199)
);

sky130_fd_sc_hd__mux4_2 c281(
.A0(net194),
.A1(in2),
.A2(net198),
.A3(net186),
.S0(in4),
.S1(net184),
.X(net200)
);

sky130_fd_sc_hd__inv_1 c282(
.A(net747),
.Y(net201)
);

sky130_fd_sc_hd__mux4_1 c283(
.A0(net69),
.A1(net199),
.A2(net192),
.A3(net198),
.S0(in17),
.S1(net194),
.X(net202)
);

sky130_fd_sc_hd__nor3b_4 c284(
.A(net199),
.B(net193),
.C_N(net839),
.Y(net203)
);

sky130_fd_sc_hd__mux4_4 c285(
.A0(net201),
.A1(net195),
.A2(net203),
.A3(out7),
.S0(net815),
.S1(net829),
.X(net204)
);

sky130_fd_sc_hd__inv_1 c286(
.A(net746),
.Y(net205)
);

sky130_fd_sc_hd__nand2_4 c287(
.A(in30),
.B(in34),
.Y(net206)
);

sky130_fd_sc_hd__nand2_2 c288(
.A(net203),
.B(net190),
.Y(net207)
);

sky130_fd_sc_hd__nor2_4 c289(
.A(net65),
.B(net74),
.Y(net208)
);

sky130_fd_sc_hd__inv_1 c290(
.A(net655),
.Y(net209)
);

sky130_fd_sc_hd__buf_1 c291(
.A(net781),
.X(net210)
);

sky130_fd_sc_hd__sdfbbn_1 c292(
.D(net199),
.RESET_B(net207),
.SCD(net190),
.SCE(net206),
.SET_B(net828),
.CLK_N(clk),
.Q(net212),
.Q_N(net211)
);

sky130_fd_sc_hd__clkinv_16 c293(
.A(net655),
.Y(net213)
);

sky130_fd_sc_hd__a2111o_2 c294(
.A1(net195),
.A2(net212),
.B1(out6),
.C1(net208),
.D1(net749),
.X(net214)
);

sky130_fd_sc_hd__sdfsbp_1 c295(
.D(net208),
.SCD(net775),
.SCE(net792),
.SET_B(net828),
.CLK(clk),
.Q(net216),
.Q_N(net215)
);

sky130_fd_sc_hd__clkbuf_16 c296(
.A(net728),
.X(net217)
);

sky130_fd_sc_hd__buf_4 c297(
.A(net815),
.X(net218)
);

sky130_fd_sc_hd__dlygate4sd1_1 c298(
.A(net767),
.X(net219)
);

sky130_fd_sc_hd__mux4_1 c299(
.A0(net190),
.A1(net196),
.A2(net93),
.A3(net216),
.S0(net206),
.S1(net207),
.X(net220)
);

sky130_fd_sc_hd__and3_1 c300(
.A(net85),
.B(net67),
.C(net770),
.X(net221)
);

sky130_fd_sc_hd__sdfsbp_2 c301(
.D(net217),
.SCD(net218),
.SCE(net207),
.SET_B(net208),
.CLK(clk),
.Q(net223),
.Q_N(net222)
);

sky130_fd_sc_hd__inv_16 c302(
.A(net747),
.Y(net224)
);

sky130_fd_sc_hd__sdfbbn_2 c303(
.D(net207),
.RESET_B(net224),
.SCD(net222),
.SCE(net211),
.SET_B(net103),
.CLK_N(clk),
.Q(out9),
.Q_N(net225)
);

sky130_fd_sc_hd__or4bb_4 c304(
.A(net224),
.B(net223),
.C_N(in25),
.D_N(net770),
.X(net226)
);

sky130_fd_sc_hd__buf_12 c305(
.A(net781),
.X(net227)
);

sky130_fd_sc_hd__mux4_4 c306(
.A0(net227),
.A1(net222),
.A2(net215),
.A3(net201),
.S0(net225),
.S1(net792),
.X(net228)
);

sky130_fd_sc_hd__mux4_2 c307(
.A0(net212),
.A1(net227),
.A2(net217),
.A3(net207),
.S0(net206),
.S1(net228),
.X(net229)
);

sky130_fd_sc_hd__and2_1 c308(
.A(net201),
.B(in18),
.X(net230)
);

sky130_fd_sc_hd__inv_2 c309(
.A(net771),
.Y(net231)
);

sky130_fd_sc_hd__or4bb_2 c310(
.A(in50),
.B(net216),
.C_N(in43),
.D_N(net101),
.X(net232)
);

sky130_fd_sc_hd__nor2_4 c311(
.A(net3),
.B(net84),
.Y(net233)
);

sky130_fd_sc_hd__or2b_4 c312(
.A(net231),
.B_N(out9),
.X(net234)
);

sky130_fd_sc_hd__or4bb_4 c313(
.A(net117),
.B(net108),
.C_N(net101),
.D_N(net234),
.X(net235)
);

sky130_fd_sc_hd__a2111oi_2 c314(
.A1(in48),
.A2(net215),
.B1(net120),
.C1(net829),
.D1(net835),
.Y(net236)
);

sky130_fd_sc_hd__or2_2 c315(
.A(net67),
.B(net230),
.X(net237)
);

sky130_fd_sc_hd__or4bb_4 c316(
.A(net232),
.B(net230),
.C_N(net231),
.D_N(in34),
.X(net238)
);

sky130_fd_sc_hd__clkbuf_1 c317(
.A(net769),
.X(net239)
);

sky130_fd_sc_hd__buf_6 c318(
.A(net769),
.X(net240)
);

sky130_fd_sc_hd__clkbuf_16 c319(
.A(net766),
.X(net241)
);

sky130_fd_sc_hd__o2111a_2 c320(
.A1(net110),
.A2(net239),
.B1(net238),
.C1(net227),
.D1(net237),
.X(net242)
);

sky130_fd_sc_hd__mux4_4 c321(
.A0(net218),
.A1(net230),
.A2(net201),
.A3(net239),
.S0(net830),
.S1(net839),
.X(out8)
);

sky130_fd_sc_hd__inv_2 c322(
.A(net771),
.Y(out28)
);

sky130_fd_sc_hd__nor2_1 c323(
.A(net241),
.B(out28),
.Y(net243)
);

sky130_fd_sc_hd__clkinv_8 c324(
.A(net896),
.Y(net244)
);

sky130_fd_sc_hd__and3_2 c325(
.A(net243),
.B(net244),
.C(out28),
.X(net245)
);

sky130_fd_sc_hd__mux4_4 c326(
.A0(net239),
.A1(net245),
.A2(net243),
.A3(net221),
.S0(in50),
.S1(net727),
.X(net246)
);

sky130_fd_sc_hd__mux4_2 c327(
.A0(net245),
.A1(net238),
.A2(net239),
.A3(net230),
.S0(out28),
.S1(net840),
.X(net247)
);

sky130_fd_sc_hd__mux4_1 c328(
.A0(net244),
.A1(net114),
.A2(net239),
.A3(net727),
.S0(net835),
.S1(net840),
.X(net248)
);

sky130_fd_sc_hd__o2111ai_2 c329(
.A1(net239),
.A2(net241),
.B1(net234),
.C1(out28),
.D1(net727),
.Y(net249)
);

sky130_fd_sc_hd__or4bb_4 c330(
.A(in11),
.B(net234),
.C_N(net834),
.D_N(net839),
.X(net250)
);

sky130_fd_sc_hd__or4bb_2 c331(
.A(net189),
.B(net138),
.C_N(net250),
.D_N(net840),
.X(net251)
);

sky130_fd_sc_hd__nand3_4 c332(
.A(in45),
.B(net142),
.C(net131),
.Y(net252)
);

sky130_fd_sc_hd__mux4_4 c333(
.A0(net130),
.A1(net234),
.A2(net250),
.A3(in45),
.S0(out7),
.S1(out28),
.X(net253)
);

sky130_fd_sc_hd__sdfbbp_1 c334(
.D(net228),
.RESET_B(in34),
.SCD(net23),
.SCE(out28),
.SET_B(net14),
.CLK(clk),
.Q(net255),
.Q_N(net254)
);

sky130_fd_sc_hd__buf_2 c335(
.A(net724),
.X(net256)
);

sky130_fd_sc_hd__or4bb_2 c336(
.A(net132),
.B(out28),
.C_N(in61),
.D_N(net215),
.X(net257)
);

sky130_fd_sc_hd__mux4_2 c337(
.A0(net16),
.A1(net256),
.A2(net254),
.A3(net250),
.S0(net131),
.S1(net841),
.X(net258)
);

sky130_fd_sc_hd__o2111ai_4 c338(
.A1(net251),
.A2(net258),
.B1(net257),
.C1(net131),
.D1(out28),
.Y(net259)
);

sky130_fd_sc_hd__o2111ai_1 c339(
.A1(in45),
.A2(net256),
.B1(net258),
.C1(net234),
.D1(net835),
.Y(net260)
);

sky130_fd_sc_hd__nand3_2 c340(
.A(net184),
.B(net252),
.C(net841),
.Y(net261)
);

sky130_fd_sc_hd__or3_2 c341(
.A(net189),
.B(net138),
.C(net234),
.X(net262)
);

sky130_fd_sc_hd__sdfbbn_1 c342(
.D(net255),
.RESET_B(net262),
.SCD(net234),
.SCE(net793),
.SET_B(net839),
.CLK_N(clk),
.Q(net264),
.Q_N(net263)
);

sky130_fd_sc_hd__sdfstp_1 c343(
.D(net131),
.SCD(net144),
.SCE(net262),
.SET_B(net16),
.CLK(clk),
.Q(net265)
);

sky130_fd_sc_hd__sdfstp_2 c344(
.D(net262),
.SCD(out28),
.SCE(net265),
.SET_B(net840),
.CLK(clk),
.Q(net266)
);

sky130_fd_sc_hd__mux4_1 c345(
.A0(net144),
.A1(net265),
.A2(net266),
.A3(in34),
.S0(net793),
.S1(net840),
.X(net267)
);

sky130_fd_sc_hd__a2111o_2 c346(
.A1(net265),
.A2(in61),
.B1(net267),
.C1(net263),
.D1(net266),
.X(net268)
);

sky130_fd_sc_hd__mux4_4 c347(
.A0(net268),
.A1(net254),
.A2(net252),
.A3(net266),
.S0(net262),
.S1(net829),
.X(net269)
);

sky130_fd_sc_hd__mux4_4 c348(
.A0(net255),
.A1(net187),
.A2(net266),
.A3(out47),
.S0(net265),
.S1(net793),
.X(net270)
);

sky130_fd_sc_hd__mux4_4 c349(
.A0(net261),
.A1(net265),
.A2(net233),
.A3(net132),
.S0(net266),
.S1(net108),
.X(net271)
);

sky130_fd_sc_hd__mux4_2 c350(
.A0(net267),
.A1(net228),
.A2(net262),
.A3(net843),
.S0(net844),
.S1(net845),
.X(net272)
);

sky130_fd_sc_hd__mux4_1 c351(
.A0(net258),
.A1(net265),
.A2(net261),
.A3(net793),
.S0(net844),
.S1(net845),
.X(net273)
);

sky130_fd_sc_hd__or4bb_4 c352(
.A(net152),
.B(net266),
.C_N(net234),
.D_N(net793),
.X(net274)
);

sky130_fd_sc_hd__or4bb_1 c353(
.A(net148),
.B(net155),
.C_N(in18),
.D_N(net839),
.X(net275)
);

sky130_fd_sc_hd__nor3b_2 c354(
.A(net274),
.B(net105),
.C_N(net831),
.Y(out60)
);

sky130_fd_sc_hd__a2111o_4 c355(
.A1(net108),
.A2(net204),
.B1(net155),
.C1(net275),
.D1(net839),
.X(net276)
);

sky130_fd_sc_hd__sdfbbn_2 c356(
.D(in61),
.RESET_B(out60),
.SCD(net153),
.SCE(net108),
.SET_B(net275),
.CLK_N(clk),
.Q(net278),
.Q_N(net277)
);

sky130_fd_sc_hd__o2111a_2 c357(
.A1(net148),
.A2(out28),
.B1(out7),
.C1(out48),
.D1(net842),
.X(net279)
);

sky130_fd_sc_hd__o2111ai_1 c358(
.A1(net151),
.A2(out46),
.B1(net225),
.C1(net158),
.D1(net751),
.Y(net280)
);

sky130_fd_sc_hd__nand3_2 c359(
.A(net108),
.B(net825),
.C(net831),
.Y(net281)
);

sky130_fd_sc_hd__sdfstp_4 c360(
.D(net281),
.SCD(in47),
.SCE(net277),
.SET_B(net86),
.CLK(clk),
.Q(net282)
);

sky130_fd_sc_hd__mux4_4 c361(
.A0(in34),
.A1(net108),
.A2(net234),
.A3(net274),
.S0(in48),
.S1(net751),
.X(out56)
);

sky130_fd_sc_hd__a2111o_2 c362(
.A1(net153),
.A2(net257),
.B1(net148),
.C1(net155),
.D1(net839),
.X(net283)
);

sky130_fd_sc_hd__buf_1 c363(
.A(net798),
.X(net284)
);

sky130_fd_sc_hd__o2111ai_2 c364(
.A1(net280),
.A2(out60),
.B1(net148),
.C1(net275),
.D1(out21),
.Y(net285)
);

sky130_fd_sc_hd__mux4_2 c365(
.A0(net283),
.A1(net263),
.A2(net282),
.A3(net155),
.S0(net158),
.S1(out48),
.X(net286)
);

sky130_fd_sc_hd__a2111oi_4 c366(
.A1(net93),
.A2(net155),
.B1(net283),
.C1(net831),
.D1(net847),
.Y(net287)
);

sky130_fd_sc_hd__a2111oi_0 c367(
.A1(net279),
.A2(net264),
.B1(net148),
.C1(net283),
.D1(net211),
.Y(net288)
);

sky130_fd_sc_hd__or4bb_4 c368(
.A(net281),
.B(net282),
.C_N(net772),
.D_N(net792),
.X(net289)
);

sky130_fd_sc_hd__sdfbbp_1 c369(
.D(net266),
.RESET_B(net283),
.SCD(net279),
.SCE(net264),
.SET_B(net847),
.CLK(clk),
.Q(net291),
.Q_N(net290)
);

sky130_fd_sc_hd__sdfbbn_1 c370(
.D(net152),
.RESET_B(net279),
.SCD(net283),
.SCE(net148),
.SET_B(net792),
.CLK_N(clk),
.Q(net293),
.Q_N(net292)
);

sky130_fd_sc_hd__o2111a_4 c371(
.A1(out12),
.A2(out23),
.B1(net292),
.C1(net772),
.D1(net792),
.X(net294)
);

sky130_fd_sc_hd__sdfbbn_2 c372(
.D(net294),
.RESET_B(net280),
.SCD(net274),
.SCE(net279),
.SET_B(out48),
.CLK_N(clk),
.Q(out11),
.Q_N(net295)
);

sky130_fd_sc_hd__mux4_1 c373(
.A0(net158),
.A1(net151),
.A2(net282),
.A3(out11),
.S0(net148),
.S1(net294),
.X(net296)
);

sky130_fd_sc_hd__mux4_1 c392(
.A0(out26),
.A1(out4),
.A2(out46),
.A3(out36),
.S0(out49),
.S1(net825),
.X(out32)
);

sky130_fd_sc_hd__mux4_4 c393(
.A0(net175),
.A1(out5),
.A2(out8),
.A3(out32),
.S0(out56),
.S1(net839),
.X(net297)
);

sky130_fd_sc_hd__mux4_2 c394(
.A0(net234),
.A1(net204),
.A2(out22),
.A3(out51),
.S0(out48),
.S1(out21),
.X(net298)
);

sky130_fd_sc_hd__mux4_4 c395(
.A0(out32),
.A1(out47),
.A2(net295),
.A3(out34),
.S0(out45),
.S1(net793),
.X(net299)
);

sky130_fd_sc_hd__nor2b_4 c396(
.A(net203),
.B_N(in9),
.Y(net300)
);

sky130_fd_sc_hd__inv_8 c397(
.A(net767),
.Y(net301)
);

sky130_fd_sc_hd__or2_1 c398(
.A(net182),
.B(in21),
.X(net302)
);

sky130_fd_sc_hd__dlygate4sd1_1 c399(
.A(net767),
.X(net303)
);

sky130_fd_sc_hd__nand2_1 c400(
.A(net303),
.B(net838),
.Y(net304)
);

sky130_fd_sc_hd__nand3_1 c401(
.A(in21),
.B(net67),
.C(net302),
.Y(net305)
);

sky130_fd_sc_hd__nand2_2 c402(
.A(net305),
.B(out7),
.Y(net306)
);

sky130_fd_sc_hd__inv_16 c403(
.A(net736),
.Y(net307)
);

sky130_fd_sc_hd__nand2_1 c404(
.A(net76),
.B(out7),
.Y(net308)
);

sky130_fd_sc_hd__nor3_4 c405(
.A(in2),
.B(net303),
.C(out7),
.Y(net309)
);

sky130_fd_sc_hd__or2b_1 c406(
.A(net304),
.B_N(net303),
.X(net310)
);

sky130_fd_sc_hd__or4bb_4 c407(
.A(net307),
.B(net300),
.C_N(net308),
.D_N(net310),
.X(net311)
);

sky130_fd_sc_hd__inv_16 c408(
.A(net782),
.Y(net312)
);

sky130_fd_sc_hd__nand3b_4 c409(
.A_N(net185),
.B(net312),
.C(net310),
.Y(net313)
);

sky130_fd_sc_hd__buf_4 c410(
.A(net669),
.X(net314)
);

sky130_fd_sc_hd__mux4_2 c411(
.A0(net307),
.A1(net308),
.A2(net312),
.A3(in2),
.S0(net302),
.S1(net310),
.X(net315)
);

sky130_fd_sc_hd__sedfxbp_1 c412(
.D(net301),
.DE(net306),
.SCD(net313),
.SCE(net310),
.CLK(clk),
.Q(net317),
.Q_N(net316)
);

sky130_fd_sc_hd__a2111oi_1 c413(
.A1(in11),
.A2(net314),
.B1(net316),
.C1(net304),
.D1(net310),
.Y(net318)
);

sky130_fd_sc_hd__sdfbbp_1 c414(
.D(net317),
.RESET_B(net318),
.SCD(net310),
.SCE(out7),
.SET_B(net706),
.CLK(clk),
.Q(net320),
.Q_N(net319)
);

sky130_fd_sc_hd__mux4_1 c415(
.A0(net192),
.A1(net318),
.A2(net76),
.A3(net313),
.S0(net309),
.S1(net310),
.X(net321)
);

sky130_fd_sc_hd__sedfxbp_2 c416(
.D(net188),
.DE(net316),
.SCD(net310),
.SCE(net794),
.CLK(clk),
.Q(net323),
.Q_N(net322)
);

sky130_fd_sc_hd__sedfxtp_1 c417(
.D(net313),
.DE(net316),
.SCD(net310),
.SCE(net794),
.CLK(clk),
.Q(net324)
);

sky130_fd_sc_hd__clkbuf_4 c418(
.A(net802),
.X(net325)
);

sky130_fd_sc_hd__and3b_2 c419(
.A_N(net324),
.B(net322),
.C(net749),
.X(net326)
);

sky130_fd_sc_hd__buf_4 c420(
.A(net802),
.X(out16)
);

sky130_fd_sc_hd__and3b_2 c421(
.A_N(net67),
.B(out16),
.C(net226),
.X(net327)
);

sky130_fd_sc_hd__mux4_1 c422(
.A0(net314),
.A1(net325),
.A2(net318),
.A3(net303),
.S0(net326),
.S1(net226),
.X(net328)
);

sky130_fd_sc_hd__or4bb_4 c423(
.A(net103),
.B(net327),
.C_N(net319),
.D_N(net310),
.X(net329)
);

sky130_fd_sc_hd__buf_6 c424(
.A(net773),
.X(net330)
);

sky130_fd_sc_hd__buf_12 c425(
.A(net896),
.X(net331)
);

sky130_fd_sc_hd__clkbuf_2 c426(
.A(net813),
.X(net332)
);

sky130_fd_sc_hd__a2111oi_2 c427(
.A1(net213),
.A2(net85),
.B1(net223),
.C1(net330),
.D1(net310),
.Y(net333)
);

sky130_fd_sc_hd__clkinv_4 c428(
.A(net782),
.Y(net334)
);

sky130_fd_sc_hd__sedfxtp_2 c429(
.D(net223),
.DE(net300),
.SCD(net325),
.SCE(net213),
.CLK(clk),
.Q(net335)
);

sky130_fd_sc_hd__nand3b_4 c430(
.A_N(net326),
.B(in35),
.C(net222),
.Y(net336)
);

sky130_fd_sc_hd__or4bb_2 c431(
.A(net331),
.B(net213),
.C_N(out16),
.D_N(net310),
.X(net337)
);

sky130_fd_sc_hd__o2111a_4 c432(
.A1(net226),
.A2(net326),
.B1(net209),
.C1(net204),
.D1(net189),
.X(net338)
);

sky130_fd_sc_hd__o2111ai_4 c433(
.A1(net219),
.A2(net103),
.B1(in35),
.C1(net225),
.D1(net788),
.Y(net339)
);

sky130_fd_sc_hd__buf_8 c434(
.A(net767),
.X(net340)
);

sky130_fd_sc_hd__sdfbbn_1 c435(
.D(net336),
.RESET_B(net335),
.SCD(net337),
.SCE(net330),
.SET_B(net788),
.CLK_N(clk),
.Q(net342),
.Q_N(net341)
);

sky130_fd_sc_hd__mux4_1 c436(
.A0(net332),
.A1(net341),
.A2(net337),
.A3(net310),
.S0(out7),
.S1(net838),
.X(net343)
);

sky130_fd_sc_hd__mux4_4 c437(
.A0(net329),
.A1(net342),
.A2(net323),
.A3(net318),
.S0(net707),
.S1(net848),
.X(net344)
);

sky130_fd_sc_hd__mux4_4 c438(
.A0(net342),
.A1(net340),
.A2(net203),
.A3(net806),
.S0(net838),
.S1(net848),
.X(net345)
);

sky130_fd_sc_hd__mux4_2 c439(
.A0(net300),
.A1(net330),
.A2(net341),
.A3(net223),
.S0(net345),
.S1(net848),
.X(net346)
);

sky130_fd_sc_hd__and3_4 c440(
.A(in2),
.B(in43),
.C(net848),
.X(net347)
);

sky130_fd_sc_hd__buf_4 c441(
.A(net796),
.X(net348)
);

sky130_fd_sc_hd__and2_0 c442(
.A(net248),
.B(net347),
.X(net349)
);

sky130_fd_sc_hd__and2_1 c443(
.A(net347),
.B(net67),
.X(net350)
);

sky130_fd_sc_hd__buf_2 c444(
.A(net796),
.X(net351)
);

sky130_fd_sc_hd__nor3b_4 c445(
.A(net350),
.B(net351),
.C_N(net849),
.Y(net352)
);

sky130_fd_sc_hd__or4bb_4 c446(
.A(net114),
.B(net249),
.C_N(net350),
.D_N(net310),
.X(out13)
);

sky130_fd_sc_hd__a2111o_4 c447(
.A1(net85),
.A2(net73),
.B1(in2),
.C1(out13),
.D1(net351),
.X(net353)
);

sky130_fd_sc_hd__or4bb_2 c448(
.A(net333),
.B(net227),
.C_N(out28),
.D_N(net85),
.X(net354)
);

sky130_fd_sc_hd__sedfxtp_4 c449(
.D(net351),
.DE(net347),
.SCD(out13),
.SCE(net350),
.CLK(clk),
.Q(net355)
);

sky130_fd_sc_hd__mux4_4 c450(
.A0(out16),
.A1(net355),
.A2(net230),
.A3(out6),
.S0(out13),
.S1(net803),
.X(net356)
);

sky130_fd_sc_hd__or4bb_1 c451(
.A(net355),
.B(net351),
.C_N(in25),
.D_N(net806),
.X(net357)
);

sky130_fd_sc_hd__mux4_2 c452(
.A0(net221),
.A1(net73),
.A2(net351),
.A3(net333),
.S0(net347),
.S1(net211),
.X(net358)
);

sky130_fd_sc_hd__or4bb_1 c453(
.A(net351),
.B(net355),
.C_N(net787),
.D_N(net833),
.X(net359)
);

sky130_fd_sc_hd__sdfbbn_2 c454(
.D(net357),
.RESET_B(net355),
.SCD(net216),
.SCE(net351),
.SET_B(out13),
.CLK_N(clk),
.Q(net361),
.Q_N(net360)
);

sky130_fd_sc_hd__mux4_2 c455(
.A0(net361),
.A1(net355),
.A2(net359),
.A3(net313),
.S0(net347),
.S1(out13),
.X(net362)
);

sky130_fd_sc_hd__mux4_1 c456(
.A0(net319),
.A1(net361),
.A2(net85),
.A3(net348),
.S0(net787),
.S1(net803),
.X(net363)
);

sky130_fd_sc_hd__mux4_4 c457(
.A0(net359),
.A1(net363),
.A2(net361),
.A3(in6),
.S0(out13),
.S1(net351),
.X(net364)
);

sky130_fd_sc_hd__mux4_4 c458(
.A0(net236),
.A1(net361),
.A2(net363),
.A3(net355),
.S0(net319),
.S1(out35),
.X(net365)
);

sky130_fd_sc_hd__mux4_1 c459(
.A0(net184),
.A1(net360),
.A2(net351),
.A3(net350),
.S0(net806),
.S1(net850),
.X(net366)
);

sky130_fd_sc_hd__mux4_4 c460(
.A0(net336),
.A1(net366),
.A2(net351),
.A3(net355),
.S0(net360),
.S1(net782),
.X(net367)
);

sky130_fd_sc_hd__mux4_1 c461(
.A0(net366),
.A1(net122),
.A2(in43),
.A3(net360),
.S0(out43),
.S1(net851),
.X(net368)
);

sky130_fd_sc_hd__nand3_2 c462(
.A(net119),
.B(net263),
.C(net252),
.Y(net369)
);

sky130_fd_sc_hd__nor3b_2 c463(
.A(net25),
.B(net86),
.C_N(out28),
.Y(net370)
);

sky130_fd_sc_hd__clkbuf_4 c464(
.A(net798),
.X(net371)
);

sky130_fd_sc_hd__nand3b_4 c465(
.A_N(net256),
.B(net233),
.C(net348),
.Y(net372)
);

sky130_fd_sc_hd__buf_8 c466(
.A(net798),
.X(net373)
);

sky130_fd_sc_hd__nand2_4 c467(
.A(net23),
.B(out21),
.Y(net374)
);

sky130_fd_sc_hd__and3b_4 c468(
.A_N(net138),
.B(net310),
.C(net846),
.X(net375)
);

sky130_fd_sc_hd__nor2b_2 c469(
.A(net216),
.B_N(out28),
.Y(net376)
);

sky130_fd_sc_hd__clkbuf_8 c470(
.A(net790),
.X(net377)
);

sky130_fd_sc_hd__and3_4 c471(
.A(net371),
.B(net377),
.C(out21),
.X(out39)
);

sky130_fd_sc_hd__inv_8 c472(
.A(net795),
.Y(net378)
);

sky130_fd_sc_hd__mux4_4 c473(
.A0(net378),
.A1(net142),
.A2(net216),
.A3(net14),
.S0(out43),
.S1(net843),
.X(net379)
);

sky130_fd_sc_hd__nand2b_2 c474(
.A_N(net348),
.B(net73),
.Y(net380)
);

sky130_fd_sc_hd__mux4_2 c475(
.A0(net250),
.A1(net327),
.A2(net23),
.A3(net93),
.S0(net377),
.S1(out13),
.X(net381)
);

sky130_fd_sc_hd__buf_16 c476(
.A(net798),
.X(net382)
);

sky130_fd_sc_hd__inv_6 c477(
.A(net795),
.Y(net383)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c478(
.A(net766),
.X(net384)
);

sky130_fd_sc_hd__buf_4 c479(
.A(net766),
.X(net385)
);

sky130_fd_sc_hd__and3b_1 c480(
.A_N(net327),
.B(net384),
.C(net844),
.X(net386)
);

sky130_fd_sc_hd__clkinv_2 c481(
.A(net766),
.Y(net387)
);

sky130_fd_sc_hd__nor3_1 c482(
.A(net382),
.B(net384),
.C(net818),
.Y(net388)
);

sky130_fd_sc_hd__mux4_4 c483(
.A0(net386),
.A1(net349),
.A2(in48),
.A3(net233),
.S0(out7),
.S1(net818),
.X(net389)
);

sky130_fd_sc_hd__a2111oi_0 c484(
.A1(net29),
.A2(out28),
.B1(net290),
.C1(in48),
.D1(net845),
.Y(net390)
);

sky130_fd_sc_hd__sdfbbp_1 c485(
.D(net212),
.RESET_B(net296),
.SCD(net29),
.SCE(net295),
.SET_B(out12),
.CLK(clk),
.Q(net392),
.Q_N(net391)
);

sky130_fd_sc_hd__a2111oi_0 c486(
.A1(net291),
.A2(net296),
.B1(net212),
.C1(net844),
.D1(net845),
.Y(net393)
);

sky130_fd_sc_hd__a2111oi_0 c487(
.A1(net385),
.A2(net390),
.B1(net275),
.C1(net376),
.D1(out28),
.Y(net394)
);

sky130_fd_sc_hd__a2111o_2 c488(
.A1(net392),
.A2(out12),
.B1(out15),
.C1(out28),
.D1(out37),
.X(net395)
);

sky130_fd_sc_hd__a2111oi_0 c489(
.A1(net349),
.A2(out22),
.B1(out6),
.C1(net395),
.D1(net376),
.Y(net396)
);

sky130_fd_sc_hd__mux4_4 c490(
.A0(net31),
.A1(net277),
.A2(net284),
.A3(out12),
.S0(out40),
.S1(net818),
.X(net397)
);

sky130_fd_sc_hd__mux4_1 c491(
.A0(net278),
.A1(net310),
.A2(out15),
.A3(net14),
.S0(net275),
.S1(net395),
.X(net398)
);

sky130_fd_sc_hd__a2111o_2 c492(
.A1(net395),
.A2(net391),
.B1(net397),
.C1(net46),
.D1(out37),
.X(net399)
);

sky130_fd_sc_hd__sdfbbn_1 c493(
.D(net291),
.RESET_B(out15),
.SCD(net275),
.SCE(in48),
.SET_B(net204),
.CLK_N(clk),
.Q(out42),
.Q_N(net400)
);

sky130_fd_sc_hd__mux4_1 c494(
.A0(net296),
.A1(net384),
.A2(out41),
.A3(net832),
.S0(net842),
.S1(net847),
.X(net401)
);

sky130_fd_sc_hd__mux4_1 c495(
.A0(net390),
.A1(out23),
.A2(net384),
.A3(net400),
.S0(net29),
.S1(net395),
.X(net402)
);

sky130_fd_sc_hd__a2111oi_2 c496(
.A1(net390),
.A2(net400),
.B1(out12),
.C1(in48),
.D1(out33),
.Y(out31)
);

sky130_fd_sc_hd__sdfbbn_2 c497(
.D(net105),
.RESET_B(out31),
.SCD(net14),
.SCE(out42),
.SET_B(net376),
.CLK_N(clk),
.Q(net404),
.Q_N(net403)
);

sky130_fd_sc_hd__a2111oi_1 c498(
.A1(net395),
.A2(net404),
.B1(net284),
.C1(net42),
.D1(net829),
.Y(out27)
);

sky130_fd_sc_hd__o2111a_2 c499(
.A1(net402),
.A2(net290),
.B1(in48),
.C1(out41),
.D1(net844),
.X(net405)
);

sky130_fd_sc_hd__o2111a_2 c500(
.A1(net31),
.A2(net404),
.B1(net395),
.C1(net391),
.D1(out37),
.X(net406)
);

sky130_fd_sc_hd__mux4_2 c501(
.A0(net264),
.A1(net284),
.A2(net278),
.A3(net397),
.S0(in48),
.S1(out41),
.X(net407)
);

sky130_fd_sc_hd__sdfbbp_1 c502(
.D(net388),
.RESET_B(out23),
.SCD(net406),
.SCE(net5),
.SET_B(net824),
.CLK(clk),
.Q(out17),
.Q_N(net408)
);

sky130_fd_sc_hd__mux4_2 c503(
.A0(net406),
.A1(net403),
.A2(net46),
.A3(net397),
.S0(out8),
.S1(net783),
.X(net409)
);

sky130_fd_sc_hd__mux4_4 c504(
.A0(net404),
.A1(in48),
.A2(net310),
.A3(in25),
.S0(out15),
.S1(net406),
.X(net410)
);

sky130_fd_sc_hd__mux4_1 c505(
.A0(net384),
.A1(net406),
.A2(net403),
.A3(net408),
.S0(net42),
.S1(out24),
.X(net411)
);

sky130_fd_sc_hd__and2_4 c528(
.A(net75),
.B(net193),
.X(net412)
);

sky130_fd_sc_hd__or2_4 c529(
.A(in4),
.B(out7),
.X(net413)
);

sky130_fd_sc_hd__nor2b_1 c530(
.A(net184),
.B_N(net826),
.Y(net414)
);

sky130_fd_sc_hd__nor2b_1 c531(
.A(net305),
.B_N(net193),
.Y(net415)
);

sky130_fd_sc_hd__inv_6 c532(
.A(net651),
.Y(net416)
);

sky130_fd_sc_hd__dlygate4sd1_1 c533(
.A(net651),
.X(net417)
);

sky130_fd_sc_hd__or2_4 c534(
.A(in17),
.B(in4),
.X(net418)
);

sky130_fd_sc_hd__inv_1 c535(
.A(net714),
.Y(net419)
);

sky130_fd_sc_hd__nand2_2 c536(
.A(net418),
.B(net312),
.Y(net420)
);

sky130_fd_sc_hd__and2_0 c537(
.A(net420),
.B(net418),
.X(net421)
);

sky130_fd_sc_hd__a2111o_4 c538(
.A1(net412),
.A2(net414),
.B1(net318),
.C1(net413),
.D1(in9),
.X(net422)
);

sky130_fd_sc_hd__clkbuf_1 c539(
.A(net736),
.X(net423)
);

sky130_fd_sc_hd__inv_1 c540(
.A(net800),
.Y(net424)
);

sky130_fd_sc_hd__buf_6 c541(
.A(net800),
.X(net425)
);

sky130_fd_sc_hd__nor2_4 c542(
.A(net302),
.B(net420),
.Y(net426)
);

sky130_fd_sc_hd__inv_4 c543(
.A(net669),
.Y(net427)
);

sky130_fd_sc_hd__nor2b_4 c544(
.A(net425),
.B_N(net416),
.Y(net428)
);

sky130_fd_sc_hd__mux4_2 c545(
.A0(net302),
.A1(net426),
.A2(net413),
.A3(net414),
.S0(net415),
.S1(net737),
.X(net429)
);

sky130_fd_sc_hd__and2_2 c546(
.A(net423),
.B(net418),
.X(net430)
);

sky130_fd_sc_hd__mux4_2 c547(
.A0(net204),
.A1(net184),
.A2(net430),
.A3(in9),
.S0(net415),
.S1(net737),
.X(net431)
);

sky130_fd_sc_hd__and2_1 c548(
.A(net430),
.B(net420),
.X(net432)
);

sky130_fd_sc_hd__mux4_2 c549(
.A0(net419),
.A1(net432),
.A2(net71),
.A3(net420),
.S0(net430),
.S1(net855),
.X(net433)
);

sky130_fd_sc_hd__clkbuf_2 c550(
.A(net784),
.X(net434)
);

sky130_fd_sc_hd__and3_1 c551(
.A(net325),
.B(net806),
.C(net857),
.X(net435)
);

sky130_fd_sc_hd__buf_4 c552(
.A(net784),
.X(net436)
);

sky130_fd_sc_hd__nand3b_1 c553(
.A_N(net86),
.B(net855),
.C(net856),
.Y(net437)
);

sky130_fd_sc_hd__or4bb_1 c554(
.A(net100),
.B(net414),
.C_N(net330),
.D_N(net310),
.X(net438)
);

sky130_fd_sc_hd__sdfrbp_1 c555(
.D(net318),
.RESET_B(net435),
.SCD(net854),
.SCE(net856),
.CLK(clk),
.Q(net440),
.Q_N(net439)
);

sky130_fd_sc_hd__or4bb_2 c556(
.A(net325),
.B(net435),
.C_N(net335),
.D_N(net332),
.X(net441)
);

sky130_fd_sc_hd__nor3_4 c557(
.A(net205),
.B(net436),
.C(net704),
.Y(net442)
);

sky130_fd_sc_hd__buf_1 c558(
.A(net797),
.X(net443)
);

sky130_fd_sc_hd__sdfrbp_2 c559(
.D(net335),
.RESET_B(net414),
.SCD(net318),
.SCE(net227),
.CLK(clk),
.Q(net445),
.Q_N(net444)
);

sky130_fd_sc_hd__mux4_2 c560(
.A0(net435),
.A1(net445),
.A2(net442),
.A3(net437),
.S0(net441),
.S1(net434),
.X(net446)
);

sky130_fd_sc_hd__buf_16 c561(
.A(net780),
.X(net447)
);

sky130_fd_sc_hd__and3_4 c562(
.A(net441),
.B(net857),
.C(net858),
.X(net448)
);

sky130_fd_sc_hd__o2111a_4 c563(
.A1(net205),
.A2(net443),
.B1(net441),
.C1(net339),
.D1(net444),
.X(out3)
);

sky130_fd_sc_hd__mux4_2 c564(
.A0(net208),
.A1(net441),
.A2(net442),
.A3(net448),
.S0(net447),
.S1(net439),
.X(net449)
);

sky130_fd_sc_hd__inv_16 c565(
.A(net773),
.Y(net450)
);

sky130_fd_sc_hd__mux4_1 c566(
.A0(net436),
.A1(net445),
.A2(net345),
.A3(net442),
.S0(net437),
.S1(net859),
.X(net451)
);

sky130_fd_sc_hd__mux4_4 c567(
.A0(net413),
.A1(net440),
.A2(net444),
.X(net452),
.S0(net761),
.S1(net859)
);

sky130_fd_sc_hd__buf_8 c568(
.A(net814),
.X(net453)
);

sky130_fd_sc_hd__mux4_4 c569(
.A0(net441),
.A1(net453),
.A2(net318),
.A3(net345),
.S0(net704),
.S1(net858),
.X(net454)
);

sky130_fd_sc_hd__mux4_2 c570(
.A0(net447),
.A1(net206),
.A2(net453),
.A3(net445),
.S0(net756),
.S1(net848),
.X(net455)
);

sky130_fd_sc_hd__mux4_4 c571(
.A0(net435),
.A1(out3),
.A2(net453),
.A3(net455),
.S0(net756),
.S1(net858),
.X(net456)
);

sky130_fd_sc_hd__or2_4 c572(
.A(net434),
.B(net851),
.X(out19)
);

sky130_fd_sc_hd__or4bb_1 c573(
.A(net443),
.B(in25),
.C_N(net453),
.D_N(net432),
.X(net457)
);

sky130_fd_sc_hd__or4bb_4 c574(
.A(net249),
.B(net350),
.C_N(net206),
.D_N(net240),
.X(net458)
);

sky130_fd_sc_hd__nor3_2 c575(
.A(net227),
.B(net120),
.C(net855),
.Y(net459)
);

sky130_fd_sc_hd__nor2_4 c576(
.A(net459),
.B(net350),
.Y(net460)
);

sky130_fd_sc_hd__sdfrtn_1 c577(
.D(net240),
.RESET_B(net458),
.SCD(net428),
.SCE(net310),
.CLK_N(clk),
.Q(net461)
);

sky130_fd_sc_hd__sdfrtp_1 c578(
.D(net432),
.RESET_B(net310),
.SCD(net84),
.SCE(net851),
.CLK(clk),
.Q(net462)
);

sky130_fd_sc_hd__clkbuf_8 c579(
.A(net800),
.X(net463)
);

sky130_fd_sc_hd__nor2b_1 c580(
.A(net227),
.B_N(net461),
.Y(net464)
);

sky130_fd_sc_hd__sdfrtp_2 c581(
.D(net230),
.RESET_B(net464),
.SCD(net461),
.SCE(out13),
.CLK(clk),
.Q(net465)
);

sky130_fd_sc_hd__nor3_4 c582(
.A(net453),
.B(net240),
.C(net428),
.Y(net466)
);

sky130_fd_sc_hd__or4bb_4 c583(
.A(net461),
.B(net230),
.C_N(net463),
.D_N(net465),
.X(net467)
);

sky130_fd_sc_hd__sdfrtp_4 c584(
.D(net118),
.RESET_B(net461),
.SCD(net416),
.SCE(out13),
.CLK(clk),
.Q(net468)
);

sky130_fd_sc_hd__o2111ai_2 c585(
.A1(net467),
.A2(net461),
.B1(net341),
.C1(net442),
.D1(net850),
.Y(net469)
);

sky130_fd_sc_hd__buf_2 c586(
.A(net800),
.X(net470)
);

sky130_fd_sc_hd__a2111o_4 c587(
.A1(net342),
.A2(net249),
.B1(net470),
.C1(in6),
.D1(net468),
.X(net471)
);

sky130_fd_sc_hd__mux4_1 c588(
.A0(net345),
.A1(net310),
.A2(net437),
.A3(net443),
.S0(net471),
.S1(out19),
.X(net472)
);

sky130_fd_sc_hd__mux4_4 c589(
.A0(net468),
.A1(net465),
.A2(net320),
.A3(net470),
.S0(net463),
.S1(net854),
.X(net473)
);

sky130_fd_sc_hd__sdfsbp_1 c590(
.D(net350),
.SCD(net471),
.SCE(net473),
.SET_B(net794),
.CLK(clk),
.Q(net475),
.Q_N(net474)
);

sky130_fd_sc_hd__mux4_1 c591(
.A0(out3),
.A1(net473),
.A2(net475),
.A3(net470),
.S0(net206),
.S1(net792),
.X(net476)
);

sky130_fd_sc_hd__mux4_2 c592(
.A0(net471),
.A1(net466),
.A2(net475),
.A3(net455),
.S0(net473),
.S1(net465),
.X(net477)
);

sky130_fd_sc_hd__a2111o_4 c593(
.A1(net473),
.A2(net474),
.B1(net204),
.C1(net470),
.D1(net761),
.X(net478)
);

sky130_fd_sc_hd__or3_2 c594(
.A(net187),
.B(net233),
.C(net799),
.X(net479)
);

sky130_fd_sc_hd__nor3b_4 c595(
.A(net142),
.B(net470),
.C_N(net791),
.Y(net480)
);

sky130_fd_sc_hd__and3b_4 c596(
.A_N(net320),
.B(net387),
.C(net377),
.X(net481)
);

sky130_fd_sc_hd__and3_1 c597(
.A(net142),
.B(net481),
.C(net846),
.X(net482)
);

sky130_fd_sc_hd__mux4_4 c598(
.A0(net387),
.A1(net86),
.A2(net481),
.A3(net383),
.S0(net14),
.S1(net416),
.X(net483)
);

sky130_fd_sc_hd__mux4_1 c599(
.A0(net458),
.A1(net310),
.A2(out8),
.A3(net377),
.S0(net846),
.S1(net861),
.X(net484)
);

sky130_fd_sc_hd__clkinv_8 c600(
.A(net805),
.Y(net485)
);

sky130_fd_sc_hd__or4bb_1 c601(
.A(net440),
.B(net481),
.C_N(out3),
.D_N(net93),
.X(net486)
);

sky130_fd_sc_hd__mux4_2 c602(
.A0(net413),
.A1(net437),
.A2(net416),
.A3(net458),
.S0(net461),
.S1(net225),
.X(net487)
);

sky130_fd_sc_hd__or4bb_1 c603(
.A(net233),
.B(net804),
.C_N(net848),
.D_N(net861),
.X(net488)
);

sky130_fd_sc_hd__clkbuf_1 c604(
.A(net805),
.X(net489)
);

sky130_fd_sc_hd__or4bb_2 c605(
.A(net458),
.B(net812),
.C_N(net833),
.D_N(net848),
.X(net490)
);

sky130_fd_sc_hd__inv_16 c606(
.A(net797),
.Y(net491)
);

sky130_fd_sc_hd__mux4_1 c607(
.A0(net482),
.A1(net73),
.A2(net5),
.A3(out13),
.S0(net862),
.S1(net864),
.X(net492)
);

sky130_fd_sc_hd__sdfbbn_1 c608(
.D(net480),
.RESET_B(out13),
.SCD(net142),
.SCE(net377),
.SET_B(net794),
.CLK_N(clk),
.Q(net494),
.Q_N(net493)
);

sky130_fd_sc_hd__mux4_2 c609(
.A0(net491),
.A1(net184),
.A2(net493),
.A3(net809),
.S0(net861),
.S1(net863),
.X(net495)
);

sky130_fd_sc_hd__mux4_4 c610(
.A0(net485),
.A1(net413),
.A2(net142),
.A3(net463),
.S0(net782),
.S1(net846),
.X(net496)
);

sky130_fd_sc_hd__mux4_4 c611(
.A0(net494),
.A1(net488),
.A2(net785),
.A3(net809),
.S0(net848),
.S1(net863),
.X(net497)
);

sky130_fd_sc_hd__mux4_2 c612(
.A0(net383),
.A1(net481),
.A2(net493),
.A3(net846),
.S0(net864),
.S1(out10),
.X(net498)
);

sky130_fd_sc_hd__mux4_2 c613(
.A0(net498),
.A1(net494),
.A2(in18),
.A3(net413),
.S0(out13),
.S1(net862),
.X(net499)
);

sky130_fd_sc_hd__mux4_1 c614(
.A0(net488),
.A1(net498),
.A2(net493),
.A3(net785),
.S0(net862),
.S1(net865),
.X(net500)
);

sky130_fd_sc_hd__mux4_1 c615(
.A0(net494),
.A1(out8),
.A2(out21),
.A3(net864),
.S0(net865),
.S1(net866),
.X(net501)
);

sky130_fd_sc_hd__mux4_4 c616(
.A0(net282),
.A1(in25),
.A2(net437),
.A3(net833),
.S0(net847),
.S1(net852),
.X(net502)
);

sky130_fd_sc_hd__mux4_2 c617(
.A0(net416),
.A1(out9),
.A2(net397),
.A3(out13),
.S0(out8),
.S1(net856),
.X(net503)
);

sky130_fd_sc_hd__mux4_1 c618(
.A0(net282),
.A1(out8),
.A2(net824),
.A3(net843),
.S0(net856),
.S1(net867),
.X(net504)
);

sky130_fd_sc_hd__mux4_1 c619(
.A0(out17),
.A1(net86),
.A2(out16),
.A3(net376),
.S0(net799),
.S1(net865),
.X(net505)
);

sky130_fd_sc_hd__mux4_4 c620(
.A0(net437),
.A1(net293),
.A2(out17),
.A3(net824),
.S0(net843),
.S1(net867),
.X(net506)
);

sky130_fd_sc_hd__mux4_1 c621(
.A0(net14),
.A1(net5),
.A2(net377),
.A3(out12),
.S0(net284),
.S1(net408),
.X(net507)
);

sky130_fd_sc_hd__mux4_4 c622(
.A0(out13),
.A1(net376),
.A2(net14),
.A3(net824),
.S0(net843),
.S1(net858),
.X(net508)
);

sky130_fd_sc_hd__mux4_4 c623(
.A0(net397),
.A1(out8),
.A2(net275),
.A3(net437),
.S0(out15),
.S1(net784),
.X(net509)
);

sky130_fd_sc_hd__mux4_4 c624(
.A0(net5),
.A1(net14),
.A2(out13),
.A3(out15),
.S0(net204),
.S1(net847),
.X(net510)
);

sky130_fd_sc_hd__mux4_4 c625(
.A0(net257),
.A1(net284),
.A2(out13),
.A3(in25),
.S0(net474),
.S1(net865),
.X(net511)
);

sky130_fd_sc_hd__mux4_4 c626(
.A0(net504),
.A1(net437),
.A2(out8),
.A3(out17),
.S0(net5),
.S1(out10),
.X(net512)
);

sky130_fd_sc_hd__o2111ai_1 c627(
.A1(net282),
.A2(out7),
.B1(net783),
.C1(out2),
.D1(net868),
.Y(net513)
);

sky130_fd_sc_hd__mux4_1 c628(
.A0(net392),
.A1(net86),
.A2(net93),
.A3(out15),
.S0(out20),
.S1(net868),
.X(out18)
);

sky130_fd_sc_hd__mux4_4 c629(
.A0(net121),
.A1(net392),
.A2(out8),
.A3(net397),
.S0(net783),
.S1(net868),
.X(net514)
);

sky130_fd_sc_hd__mux4_1 c630(
.A0(net392),
.A1(net505),
.A2(out18),
.A3(net310),
.S0(net833),
.S1(out10),
.X(net515)
);

sky130_fd_sc_hd__mux4_1 c631(
.A0(out9),
.A1(net397),
.A2(net408),
.A3(net810),
.S0(net867),
.S1(net868),
.X(net516)
);

sky130_fd_sc_hd__mux4_4 c632(
.A0(out13),
.A1(net391),
.A2(net811),
.A3(net824),
.S0(out20),
.S1(net868),
.X(net517)
);

sky130_fd_sc_hd__mux4_1 c633(
.A0(net442),
.A1(net501),
.A2(out9),
.A3(net86),
.S0(net852),
.S1(net868),
.X(net518)
);

sky130_fd_sc_hd__mux4_2 c634(
.A0(net86),
.A1(net783),
.A2(net808),
.A3(net824),
.S0(net852),
.S1(net868),
.X(net519)
);

sky130_fd_sc_hd__mux4_4 c635(
.A0(net275),
.A1(net519),
.A2(out8),
.A3(net808),
.S0(net829),
.S1(net868),
.X(net520)
);

sky130_fd_sc_hd__mux4_1 c636(
.A0(net513),
.A1(net519),
.A2(net391),
.A3(net791),
.S0(net810),
.S1(net853),
.X(net521)
);

sky130_fd_sc_hd__mux4_2 c637(
.A0(net204),
.A1(net789),
.A2(net801),
.A3(net811),
.S0(net853),
.S1(out20),
.X(net522)
);

sky130_fd_sc_hd__inv_4 c660(
.A(net638),
.Y(net523)
);

sky130_fd_sc_hd__inv_16 c661(
.A(net638),
.Y(net524)
);

sky130_fd_sc_hd__clkinv_16 c662(
.A(net714),
.Y(net525)
);

sky130_fd_sc_hd__nor2_1 c663(
.A(net317),
.B(in9),
.Y(net526)
);

sky130_fd_sc_hd__and2_2 c664(
.A(net184),
.B(net427),
.X(net527)
);

sky130_fd_sc_hd__nor2_1 c665(
.A(net71),
.B(net524),
.Y(net528)
);

sky130_fd_sc_hd__nor2b_2 c666(
.A(net528),
.B_N(net424),
.Y(net529)
);

sky130_fd_sc_hd__and2b_2 c667(
.A_N(net528),
.B(net524),
.X(net530)
);

sky130_fd_sc_hd__buf_16 c668(
.A(net714),
.X(net531)
);

sky130_fd_sc_hd__and2_0 c669(
.A(net323),
.B(net424),
.X(net532)
);

sky130_fd_sc_hd__buf_12 c670(
.A(out2),
.X(net533)
);

sky130_fd_sc_hd__buf_12 c671(
.A(net714),
.X(net534)
);

sky130_fd_sc_hd__mux4_4 c672(
.A0(net427),
.A1(net529),
.A2(net531),
.A3(net323),
.S0(net524),
.S1(net193),
.X(net535)
);

sky130_fd_sc_hd__and2b_1 c673(
.A_N(net525),
.B(net872),
.X(net536)
);

sky130_fd_sc_hd__nor3b_1 c674(
.A(net531),
.B(net193),
.C_N(net871),
.Y(net537)
);

sky130_fd_sc_hd__or3b_4 c675(
.A(net536),
.B(net534),
.C_N(net872),
.X(net538)
);

sky130_fd_sc_hd__a2111oi_1 c676(
.A1(net538),
.A2(net320),
.B1(net317),
.C1(net533),
.D1(net526),
.Y(net539)
);

sky130_fd_sc_hd__dlygate4sd3_1 c677(
.A(net807),
.X(net540)
);

sky130_fd_sc_hd__sdfbbn_2 c678(
.D(net534),
.RESET_B(net532),
.SCD(net196),
.SCE(net540),
.SET_B(net871),
.CLK_N(clk),
.Q(net542),
.Q_N(net541)
);

sky130_fd_sc_hd__clkinv_8 c679(
.A(net897),
.Y(net543)
);

sky130_fd_sc_hd__mux4_4 c680(
.A0(net523),
.A1(net540),
.A2(net543),
.A3(net531),
.S0(net541),
.S1(net532),
.X(net544)
);

sky130_fd_sc_hd__o2111ai_1 c681(
.A1(net544),
.A2(net538),
.B1(net542),
.C1(net184),
.D1(net524),
.Y(net545)
);

sky130_fd_sc_hd__inv_8 c682(
.A(net773),
.Y(net546)
);

sky130_fd_sc_hd__and3_1 c683(
.A(net334),
.B(net303),
.C(net455),
.X(net547)
);

sky130_fd_sc_hd__or4bb_1 c684(
.A(net330),
.B(net432),
.C_N(net529),
.D_N(net860),
.X(net548)
);

sky130_fd_sc_hd__buf_1 c685(
.A(net814),
.X(net549)
);

sky130_fd_sc_hd__buf_1 c686(
.A(net807),
.X(net550)
);

sky130_fd_sc_hd__and3_4 c687(
.A(net533),
.B(net330),
.C(in9),
.X(net551)
);

sky130_fd_sc_hd__clkinv_8 c688(
.A(net773),
.Y(net552)
);

sky130_fd_sc_hd__inv_4 c689(
.A(net761),
.Y(net553)
);

sky130_fd_sc_hd__and3b_2 c690(
.A_N(net543),
.B(net546),
.C(net860),
.X(net554)
);

sky130_fd_sc_hd__buf_1 c691(
.A(net761),
.X(net555)
);

sky130_fd_sc_hd__or3b_2 c692(
.A(net555),
.B(net550),
.C_N(net444),
.X(net556)
);

sky130_fd_sc_hd__a2111oi_4 c693(
.A1(net303),
.A2(net529),
.B1(net330),
.C1(net556),
.D1(net541),
.Y(net557)
);

sky130_fd_sc_hd__sdfbbp_1 c694(
.D(net196),
.RESET_B(net537),
.SCD(net556),
.SCE(net455),
.SET_B(net552),
.CLK(clk),
.Q(net559),
.Q_N(net558)
);

sky130_fd_sc_hd__mux4_1 c695(
.A0(net559),
.A1(net552),
.A2(net532),
.A3(net554),
.S0(net332),
.S1(net556),
.X(net560)
);

sky130_fd_sc_hd__sdfbbn_1 c696(
.D(net545),
.RESET_B(net533),
.SCD(net549),
.SCE(net455),
.SET_B(net712),
.CLK_N(clk),
.Q(net562),
.Q_N(net561)
);

sky130_fd_sc_hd__mux4_4 c697(
.A0(net532),
.A1(net543),
.A2(net556),
.A3(net562),
.S0(net330),
.S1(net529),
.X(net563)
);

sky130_fd_sc_hd__mux4_4 c698(
.A0(net554),
.A1(net555),
.A2(net556),
.A3(net561),
.S0(net310),
.S1(net874),
.X(net564)
);

sky130_fd_sc_hd__mux4_4 c699(
.A0(net540),
.A1(net445),
.A2(net556),
.A3(net559),
.S0(net561),
.S1(net860),
.X(net565)
);

sky130_fd_sc_hd__mux4_4 c700(
.A0(net445),
.A1(net537),
.A2(net565),
.A3(net556),
.S0(net552),
.S1(net874),
.X(net566)
);

sky130_fd_sc_hd__mux4_2 c701(
.A0(net556),
.A1(net546),
.A2(net562),
.A3(net565),
.S0(net206),
.S1(net558),
.X(net567)
);

sky130_fd_sc_hd__mux4_1 c702(
.A0(net188),
.A1(net565),
.A2(net206),
.A3(net567),
.S0(net93),
.S1(net561),
.X(net568)
);

sky130_fd_sc_hd__mux4_2 c703(
.A0(net414),
.A1(net566),
.A2(net334),
.A3(net549),
.S0(net712),
.S1(net875),
.X(net569)
);

sky130_fd_sc_hd__sdfbbn_2 c704(
.D(net526),
.RESET_B(net455),
.SCD(net432),
.SCE(net84),
.SET_B(net462),
.CLK_N(clk),
.Q(net571),
.Q_N(net570)
);

sky130_fd_sc_hd__or4bb_1 c705(
.A(net566),
.B(net567),
.C_N(net565),
.D_N(net541),
.X(net572)
);

sky130_fd_sc_hd__sdfsbp_2 c706(
.D(net84),
.SCD(net571),
.SCE(net562),
.SET_B(net567),
.CLK(clk),
.Q(net574),
.Q_N(net573)
);

sky130_fd_sc_hd__sdfbbp_1 c707(
.D(in9),
.RESET_B(in43),
.SCD(out6),
.SCE(net542),
.SET_B(net553),
.CLK(clk),
.Q(net576),
.Q_N(net575)
);

sky130_fd_sc_hd__sdfbbn_1 c708(
.D(net574),
.RESET_B(net564),
.SCD(net432),
.SCE(net570),
.SET_B(net875),
.CLK_N(clk),
.Q(net578),
.Q_N(net577)
);

sky130_fd_sc_hd__mux4_2 c709(
.A0(net567),
.A1(net565),
.A2(net470),
.A3(net576),
.S0(net573),
.S1(net455),
.X(net579)
);

sky130_fd_sc_hd__or4bb_1 c710(
.A(net565),
.B(net470),
.C_N(in9),
.D_N(net876),
.X(net580)
);

sky130_fd_sc_hd__sdfbbn_2 c711(
.D(net562),
.RESET_B(net576),
.SCD(net573),
.SCE(net547),
.SET_B(net875),
.CLK_N(clk),
.Q(net582),
.Q_N(net581)
);

sky130_fd_sc_hd__mux4_4 c712(
.A0(net340),
.A1(net576),
.A2(net84),
.A3(net455),
.S0(net573),
.S1(net184),
.X(net583)
);

sky130_fd_sc_hd__mux4_4 c713(
.A0(net530),
.A1(net583),
.A2(net526),
.A3(net581),
.S0(net573),
.S1(net206),
.X(net584)
);

sky130_fd_sc_hd__a2111oi_0 c714(
.A1(net542),
.A2(net582),
.B1(net574),
.C1(in9),
.D1(net475),
.Y(net585)
);

sky130_fd_sc_hd__o2111a_4 c715(
.A1(net549),
.A2(net564),
.B1(net462),
.C1(net310),
.D1(net583),
.X(net586)
);

sky130_fd_sc_hd__mux4_4 c716(
.A0(net582),
.A1(net574),
.A2(net575),
.A3(net184),
.S0(in43),
.S1(net797),
.X(net587)
);

sky130_fd_sc_hd__mux4_2 c717(
.A0(net583),
.A1(net560),
.A2(in43),
.A3(net587),
.S0(out7),
.S1(net786),
.X(net588)
);

sky130_fd_sc_hd__mux4_1 c718(
.A0(net574),
.A1(net583),
.A2(net121),
.A3(net587),
.S0(out7),
.S1(net575),
.X(net589)
);

sky130_fd_sc_hd__mux4_2 c719(
.A0(net432),
.A1(net587),
.A2(net549),
.A3(net576),
.S0(net561),
.S1(net871),
.X(net590)
);

sky130_fd_sc_hd__mux4_4 c720(
.A0(net560),
.A1(net542),
.A2(net475),
.A3(net585),
.S0(net575),
.S1(net879),
.X(net591)
);

sky130_fd_sc_hd__a2111o_1 c721(
.A1(net206),
.A2(net583),
.B1(net553),
.C1(net566),
.D1(net876),
.X(net592)
);

sky130_fd_sc_hd__mux4_2 c722(
.A0(net553),
.A1(net585),
.A2(net574),
.A3(net577),
.S0(net455),
.S1(net756),
.X(net593)
);

sky130_fd_sc_hd__mux4_4 c723(
.A0(net591),
.A1(net470),
.A2(net593),
.A3(net797),
.S0(net877),
.S1(net879),
.X(net594)
);

sky130_fd_sc_hd__mux4_4 c724(
.A0(net585),
.A1(net593),
.A2(net580),
.A3(net530),
.S0(net575),
.S1(net860),
.X(net595)
);

sky130_fd_sc_hd__sdfbbp_1 c725(
.D(net591),
.RESET_B(net593),
.SCD(net786),
.SCE(net860),
.SET_B(net883),
.CLK(clk),
.Q(net597),
.Q_N(net596)
);

sky130_fd_sc_hd__a2111o_2 c726(
.A1(net320),
.A2(net455),
.B1(in18),
.C1(net866),
.D1(net878),
.X(net598)
);

sky130_fd_sc_hd__mux4_4 c727(
.A0(net122),
.A1(net598),
.A2(net547),
.A3(net866),
.S0(net876),
.S1(net881),
.X(net599)
);

sky130_fd_sc_hd__o2111ai_2 c728(
.A1(net596),
.A2(net865),
.B1(net866),
.C1(net873),
.D1(net878),
.Y(net600)
);

sky130_fd_sc_hd__mux4_4 c729(
.A0(net527),
.A1(net310),
.A2(net93),
.A3(net813),
.S0(net874),
.S1(net880),
.X(net601)
);

sky130_fd_sc_hd__mux4_2 c730(
.A0(net380),
.A1(net73),
.A2(net598),
.A3(net600),
.S0(net474),
.S1(net463),
.X(net602)
);

sky130_fd_sc_hd__o2111ai_1 c731(
.A1(in18),
.A2(net372),
.B1(net865),
.C1(net866),
.D1(net873),
.Y(net603)
);

sky130_fd_sc_hd__mux4_4 c732(
.A0(net332),
.A1(net598),
.A2(net570),
.A3(net600),
.S0(net813),
.S1(net873),
.X(net604)
);

sky130_fd_sc_hd__o2111a_1 c733(
.A1(net600),
.A2(in18),
.B1(net598),
.C1(net849),
.D1(net884),
.X(net605)
);

sky130_fd_sc_hd__mux4_1 c734(
.A0(net455),
.A1(net380),
.A2(net204),
.A3(in18),
.S0(net872),
.S1(net884),
.X(net606)
);

sky130_fd_sc_hd__mux4_4 c735(
.A0(net527),
.A1(in25),
.A2(net463),
.A3(net600),
.S0(net879),
.S1(net884),
.X(net607)
);

sky130_fd_sc_hd__mux4_4 c736(
.A0(net600),
.A1(net488),
.A2(net816),
.A3(net866),
.S0(net872),
.S1(net878),
.X(net608)
);

sky130_fd_sc_hd__mux4_4 c737(
.A0(net597),
.A1(net488),
.A2(net600),
.A3(net495),
.S0(net807),
.S1(net876),
.X(net609)
);

sky130_fd_sc_hd__mux4_2 c738(
.A0(net571),
.A1(net598),
.A2(out6),
.A3(net184),
.S0(net849),
.S1(net872),
.X(net610)
);

sky130_fd_sc_hd__mux4_4 c739(
.A0(net527),
.A1(net598),
.A2(net801),
.A3(net879),
.S0(net883),
.S1(net885),
.X(net611)
);

sky130_fd_sc_hd__mux4_2 c740(
.A0(net527),
.A1(net470),
.A2(net865),
.A3(net878),
.S0(net886),
.S1(net887),
.X(net612)
);

sky130_fd_sc_hd__mux4_4 c741(
.A0(net462),
.A1(in6),
.A2(net812),
.A3(net882),
.S0(net887),
.S1(net888),
.X(net613)
);

sky130_fd_sc_hd__mux4_4 c742(
.A0(net455),
.A1(net600),
.A2(net613),
.A3(net597),
.S0(net879),
.S1(net885),
.X(net614)
);

sky130_fd_sc_hd__mux4_2 c743(
.A0(net495),
.A1(net613),
.A2(net614),
.A3(net488),
.S0(net881),
.S1(net886),
.X(net615)
);

sky130_fd_sc_hd__mux4_1 c744(
.A0(net613),
.A1(net614),
.A2(net120),
.A3(net884),
.S0(net888),
.S1(net889),
.X(net616)
);

sky130_fd_sc_hd__mux4_4 c745(
.A0(net372),
.A1(net614),
.A2(in18),
.A3(net887),
.S0(net888),
.S1(net889),
.X(net617)
);

sky130_fd_sc_hd__mux4_4 c746(
.A0(net613),
.A1(net596),
.A2(net791),
.A3(net807),
.S0(net812),
.S1(net889),
.X(net618)
);

sky130_fd_sc_hd__mux4_1 c747(
.A0(net618),
.A1(net614),
.A2(in25),
.A3(net791),
.S0(net885),
.S1(net887),
.X(net619)
);

sky130_fd_sc_hd__mux4_1 c748(
.A0(net121),
.A1(net597),
.A2(net488),
.A3(net310),
.S0(net829),
.S1(net853),
.X(net620)
);

sky130_fd_sc_hd__mux4_2 c749(
.A0(net310),
.A1(net72),
.A2(net547),
.A3(net578),
.S0(net870),
.S1(net886),
.X(net621)
);

sky130_fd_sc_hd__mux4_1 c750(
.A0(net377),
.A1(net489),
.A2(net596),
.A3(net870),
.S0(net888),
.S1(net890),
.X(net622)
);

sky130_fd_sc_hd__mux4_4 c751(
.A0(net377),
.A1(net292),
.A2(net474),
.A3(net847),
.S0(net870),
.S1(net886),
.X(net623)
);

sky130_fd_sc_hd__mux4_4 c752(
.A0(net293),
.A1(net623),
.A2(net121),
.A3(net853),
.S0(net867),
.S1(net888),
.X(net624)
);

sky130_fd_sc_hd__a2111o_2 c753(
.A1(net488),
.A2(net597),
.B1(net292),
.C1(net817),
.D1(net870),
.X(net625)
);

sky130_fd_sc_hd__mux4_1 c754(
.A0(in25),
.A1(net784),
.A2(net789),
.A3(net867),
.S0(net886),
.S1(net888),
.X(net626)
);

sky130_fd_sc_hd__mux4_4 c755(
.A0(net397),
.A1(net580),
.A2(net623),
.A3(net463),
.S0(net93),
.S1(net869),
.X(net627)
);

sky130_fd_sc_hd__mux4_4 c756(
.A0(net597),
.A1(net626),
.A2(net293),
.A3(net869),
.S0(net877),
.S1(net892),
.X(net628)
);

sky130_fd_sc_hd__mux4_2 c757(
.A0(net475),
.A1(net622),
.A2(net488),
.A3(net120),
.S0(net867),
.S1(net891),
.X(net629)
);

sky130_fd_sc_hd__mux4_4 c758(
.A0(net376),
.A1(net463),
.A2(net628),
.A3(net817),
.S0(net890),
.S1(net894),
.X(net630)
);

sky130_fd_sc_hd__mux4_4 c759(
.A0(net121),
.A1(net630),
.A2(net628),
.A3(net488),
.S0(net865),
.S1(net893),
.X(net631)
);

sky130_fd_sc_hd__mux4_4 c760(
.A0(net578),
.A1(net376),
.A2(net204),
.A3(net816),
.S0(net865),
.S1(net893),
.X(net632)
);

sky130_fd_sc_hd__mux4_2 c761(
.A0(net547),
.A1(net377),
.A2(net799),
.A3(net805),
.S0(net890),
.S1(net895),
.X(net633)
);

sky130_fd_sc_hd__mux4_2 c762(
.A0(net489),
.A1(net596),
.A2(net799),
.A3(net869),
.S0(net891),
.S1(net895),
.X(net634)
);

sky130_fd_sc_hd__mux4_2 c763(
.A0(net634),
.A1(net628),
.A2(net756),
.A3(net805),
.S0(net852),
.S1(net891),
.X(net635)
);

sky130_fd_sc_hd__mux4_4 c764(
.A0(net624),
.A1(net635),
.A2(net310),
.A3(net867),
.S0(net877),
.S1(net888),
.X(net636)
);

sky130_fd_sc_hd__or4bb_4 merge765(
.A(net163),
.B(net5),
.C_N(net57),
.D_N(net176),
.X(net637)
);

sky130_fd_sc_hd__dlygate4sd3_1 merge766(
.A(net897),
.X(net638)
);

sky130_fd_sc_hd__or4bb_2 merge767(
.A(net90),
.B(in45),
.C_N(net238),
.D_N(net727),
.X(net639)
);

sky130_fd_sc_hd__or4bb_4 merge768(
.A(in59),
.B(net12),
.C_N(net30),
.D_N(in20),
.X(net640)
);

sky130_fd_sc_hd__or4bb_4 merge769(
.A(net186),
.B(net203),
.C_N(net300),
.D_N(out6),
.X(net641)
);

sky130_fd_sc_hd__mux4_4 merge770(
.A0(net18),
.A1(net225),
.A2(net437),
.A3(net479),
.S0(net482),
.S1(net804),
.X(net642)
);

sky130_fd_sc_hd__o2111a_4 merge771(
.A1(net87),
.A2(net98),
.B1(net91),
.C1(net827),
.D1(net828),
.X(net643)
);

sky130_fd_sc_hd__inv_8 merge772(
.A(net778),
.Y(net644)
);

sky130_fd_sc_hd__a2111oi_2 merge773(
.A1(net550),
.A2(net529),
.B1(net537),
.C1(net196),
.D1(net860),
.Y(net645)
);

sky130_fd_sc_hd__mux4_2 merge774(
.A0(net313),
.A1(net211),
.A2(out28),
.A3(net235),
.S0(net345),
.S1(net832),
.X(net646)
);

sky130_fd_sc_hd__mux4_4 merge775(
.A0(net428),
.A1(net233),
.A2(out13),
.A3(net469),
.S0(net460),
.S1(net468),
.X(net647)
);

sky130_fd_sc_hd__or4bb_4 merge776(
.A(net71),
.B(net70),
.C_N(net73),
.D_N(net69),
.X(net648)
);

sky130_fd_sc_hd__a2111o_4 merge777(
.A1(net324),
.A2(in35),
.B1(net318),
.C1(net707),
.D1(net749),
.X(net649)
);

sky130_fd_sc_hd__a2111oi_0 merge778(
.A1(in20),
.A2(net36),
.B1(in34),
.C1(net139),
.D1(net819),
.Y(net650)
);

sky130_fd_sc_hd__buf_2 merge779(
.A(out2),
.X(net651)
);

sky130_fd_sc_hd__or4bb_4 merge780(
.A(in7),
.B(net90),
.C_N(net109),
.D_N(net830),
.X(net652)
);

sky130_fd_sc_hd__o2111a_2 merge781(
.A1(in35),
.A2(net74),
.B1(net414),
.C1(net208),
.D1(net857),
.X(net653)
);

sky130_fd_sc_hd__or4bb_4 merge782(
.A(net352),
.B(net146),
.C_N(net306),
.D_N(net375),
.X(net654)
);

sky130_fd_sc_hd__buf_8 merge783(
.A(net771),
.X(net655)
);

sky130_fd_sc_hd__inv_6 merge784(
.A(net778),
.Y(net656)
);

sky130_fd_sc_hd__or4bb_4 merge785(
.A(net64),
.B(net72),
.C_N(net69),
.D_N(out7),
.X(net657)
);

sky130_fd_sc_hd__a2111oi_2 merge786(
.A1(net109),
.A2(net116),
.B1(in33),
.C1(net128),
.D1(net8),
.Y(net658)
);

sky130_fd_sc_hd__o2111ai_2 merge787(
.A1(net235),
.A2(net237),
.B1(net84),
.C1(net238),
.D1(out7),
.Y(net659)
);

sky130_fd_sc_hd__mux4_2 merge788(
.A0(net330),
.A1(net414),
.A2(net482),
.A3(out6),
.S0(net812),
.S1(net856),
.X(net660)
);

sky130_fd_sc_hd__a2111o_2 merge789(
.A1(net111),
.A2(net113),
.B1(net107),
.C1(net251),
.D1(net131),
.X(net661)
);

sky130_fd_sc_hd__or4bb_2 merge790(
.A(net186),
.B(net183),
.C_N(net208),
.D_N(net775),
.X(net662)
);

sky130_fd_sc_hd__or4bb_4 merge791(
.A(net424),
.B(net432),
.C_N(net414),
.D_N(net706),
.X(net663)
);

sky130_fd_sc_hd__mux4_1 merge792(
.A0(net123),
.A1(net23),
.A2(net131),
.A3(in37),
.S0(net100),
.S1(net775),
.X(net664)
);

sky130_fd_sc_hd__mux4_4 merge793(
.A0(in55),
.A1(out47),
.A2(in45),
.A3(in9),
.S0(net93),
.S1(net107),
.X(net665)
);

sky130_fd_sc_hd__or4bb_4 merge794(
.A(net421),
.B(in4),
.C_N(net306),
.D_N(net192),
.X(net666)
);

sky130_fd_sc_hd__mux4_1 merge795(
.A0(net115),
.A1(net8),
.A2(net135),
.A3(in52),
.S0(net110),
.S1(net111),
.X(net667)
);

sky130_fd_sc_hd__mux4_1 merge796(
.A0(net173),
.A1(in14),
.A2(out52),
.A3(net172),
.S0(net176),
.S1(out1),
.X(net668)
);

sky130_fd_sc_hd__sdfstp_1 merge797(
.D(net308),
.SCD(net306),
.SCE(net415),
.SET_B(net204),
.CLK(clk),
.Q(net669)
);

sky130_fd_sc_hd__mux4_4 merge798(
.A0(net13),
.A1(net12),
.A2(net19),
.A3(net5),
.S0(net8),
.S1(net819),
.X(net670)
);

sky130_fd_sc_hd__a2111o_4 merge799(
.A1(net112),
.A2(in14),
.B1(net111),
.C1(net117),
.D1(net120),
.X(net671)
);

sky130_fd_sc_hd__or4bb_2 merge800(
.A(net309),
.B(net322),
.C_N(net417),
.D_N(net413),
.X(net672)
);

sky130_fd_sc_hd__or4bb_4 merge801(
.A(net193),
.B(net194),
.C_N(in16),
.D_N(net196),
.X(net673)
);

sky130_fd_sc_hd__or4bb_2 merge802(
.A(net426),
.B(net528),
.C_N(net524),
.D_N(net530),
.X(net674)
);

sky130_fd_sc_hd__mux4_1 merge803(
.A0(net448),
.A1(net335),
.A2(net209),
.A3(net322),
.S0(net300),
.S1(net859),
.X(net675)
);

sky130_fd_sc_hd__or4bb_2 merge804(
.A(net60),
.B(net49),
.C_N(net28),
.D_N(net44),
.X(net676)
);

sky130_fd_sc_hd__mux4_2 merge805(
.A0(net61),
.A1(out49),
.A2(net163),
.A3(in54),
.S0(in48),
.S1(net14),
.X(net677)
);

sky130_fd_sc_hd__mux4_4 merge806(
.A0(net12),
.A1(in57),
.A2(net9),
.A3(in33),
.S0(net30),
.S1(net820),
.X(net678)
);

sky130_fd_sc_hd__mux4_1 merge807(
.A0(net7),
.A1(net21),
.A2(net12),
.A3(net37),
.S0(net38),
.S1(out49),
.X(net679)
);

sky130_fd_sc_hd__mux4_4 merge808(
.A0(net146),
.A1(in11),
.A2(net189),
.A3(net155),
.S0(net283),
.S1(net266),
.X(net680)
);

sky130_fd_sc_hd__mux4_2 merge809(
.A0(net369),
.A1(net306),
.A2(net376),
.A3(net134),
.S0(net8),
.S1(net23),
.X(net681)
);

sky130_fd_sc_hd__mux4_4 merge810(
.A0(net370),
.A1(net376),
.A2(net204),
.A3(net252),
.S0(net377),
.S1(net352),
.X(net682)
);

sky130_fd_sc_hd__mux4_1 merge811(
.A0(net238),
.A1(net218),
.A2(net374),
.A3(out13),
.S0(net384),
.S1(net834),
.X(net683)
);

sky130_fd_sc_hd__mux4_4 merge812(
.A0(net206),
.A1(net207),
.A2(in42),
.A3(net100),
.S0(net222),
.S1(net828),
.X(net684)
);

sky130_fd_sc_hd__mux4_2 merge813(
.A0(net373),
.A1(out8),
.A2(net306),
.A3(net375),
.S0(out13),
.S1(net384),
.X(net685)
);

sky130_fd_sc_hd__mux4_1 merge814(
.A0(net325),
.A1(net329),
.A2(net234),
.A3(net238),
.S0(out28),
.S1(net838),
.X(net686)
);

sky130_fd_sc_hd__mux4_1 merge815(
.A0(net197),
.A1(net188),
.A2(net210),
.A3(net104),
.S0(net208),
.S1(net838),
.X(net687)
);

sky130_fd_sc_hd__mux4_4 merge816(
.A0(net310),
.A1(net308),
.A2(out7),
.A3(net104),
.S0(net324),
.S1(net329),
.X(net688)
);

sky130_fd_sc_hd__a2111oi_4 merge817(
.A1(net526),
.A2(net530),
.B1(net413),
.C1(net415),
.D1(net312),
.Y(net689)
);

sky130_fd_sc_hd__mux4_2 merge818(
.A0(net197),
.A1(net329),
.A2(net310),
.A3(net133),
.S0(net140),
.S1(net136),
.X(net690)
);

sky130_fd_sc_hd__mux4_4 merge819(
.A0(in41),
.A1(net38),
.A2(out49),
.A3(in38),
.S0(net10),
.S1(net710),
.X(net691)
);

sky130_fd_sc_hd__mux4_2 merge820(
.A0(net104),
.A1(net208),
.A2(net124),
.A3(net110),
.S0(net828),
.S1(net832),
.X(net692)
);

sky130_fd_sc_hd__mux4_2 merge821(
.A0(net529),
.A1(net551),
.A2(net545),
.A3(net206),
.S0(net712),
.S1(net871),
.X(net693)
);

sky130_fd_sc_hd__mux4_1 merge822(
.A0(net207),
.A1(net190),
.A2(net208),
.A3(net8),
.S0(net92),
.S1(net16),
.X(net694)
);

sky130_fd_sc_hd__mux4_4 merge823(
.A0(net187),
.A1(net186),
.A2(net182),
.A3(out7),
.S0(net100),
.S1(net857),
.X(net695)
);

sky130_fd_sc_hd__mux4_1 merge824(
.A0(net101),
.A1(in25),
.A2(out47),
.A3(net12),
.S0(net21),
.S1(net17),
.X(net696)
);

sky130_fd_sc_hd__mux4_2 merge825(
.A0(net337),
.A1(net335),
.A2(net330),
.A3(in40),
.S0(net215),
.S1(net208),
.X(net697)
);

sky130_fd_sc_hd__mux4_4 merge826(
.A0(net55),
.A1(out47),
.A2(net140),
.A3(net131),
.S0(net138),
.S1(net837),
.X(net698)
);

sky130_fd_sc_hd__a2111o_1 merge827(
.A1(net130),
.A2(net131),
.B1(net129),
.C1(net2),
.D1(net834),
.X(net699)
);

sky130_fd_sc_hd__mux4_1 merge828(
.A0(net538),
.A1(net72),
.A2(net524),
.A3(net339),
.S0(net545),
.S1(net444),
.X(net700)
);

sky130_fd_sc_hd__mux4_4 merge829(
.A0(net450),
.A1(net428),
.A2(net437),
.A3(net529),
.S0(net537),
.S1(net712),
.X(net701)
);

sky130_fd_sc_hd__mux4_4 merge830(
.A0(net539),
.A1(net540),
.A2(net426),
.A3(net427),
.S0(net193),
.S1(net871),
.X(net702)
);

sky130_fd_sc_hd__dfrbp_1 merge831(
.Q_N(net452),
.RESET_B(net438),
.CLK(clk),
.Q(net704)
);

sky130_fd_sc_hd__nor2_1 merge832(
.A(net490),
.B(net492),
.Y(net705)
);

sky130_fd_sc_hd__dfrbp_2 merge833(
.D(net311),
.RESET_B(net315),
.CLK(clk),
.Q(net707),
.Q_N(net706)
);

sky130_fd_sc_hd__and2_0 merge834(
.A(net572),
.B(net584),
.X(net708)
);

sky130_fd_sc_hd__nor2b_1 merge835(
.A(net272),
.B_N(net259),
.Y(net709)
);

sky130_fd_sc_hd__dfrtn_1 merge836(
.D(net670),
.RESET_B(net15),
.CLK_N(clk),
.Q(net710)
);

sky130_fd_sc_hd__nand2b_4 merge837(
.A_N(net299),
.B(net297),
.Y(net711)
);

sky130_fd_sc_hd__dfrtp_1 merge838(
.D(net548),
.RESET_B(net557),
.CLK(clk),
.Q(net712)
);

sky130_fd_sc_hd__and2_0 merge839(
.A(net96),
.B(net643),
.X(net713)
);

sky130_fd_sc_hd__dfrtp_2 merge840(
.D(net663),
.RESET_B(net674),
.CLK(clk),
.Q(net714)
);

sky130_fd_sc_hd__nor2b_1 merge841(
.A(net353),
.B_N(net358),
.Y(net715)
);

sky130_fd_sc_hd__nand2_1 merge842(
.A(net381),
.B(net379),
.Y(net716)
);

sky130_fd_sc_hd__nor2b_2 merge843(
.A(net393),
.B_N(net398),
.Y(net717)
);

sky130_fd_sc_hd__dfrtp_4 merge844(
.D(net41),
.RESET_B(net640),
.CLK(clk),
.Q(net718)
);

sky130_fd_sc_hd__nor2b_4 merge845(
.A(net229),
.B_N(net214),
.Y(net719)
);

sky130_fd_sc_hd__and2b_1 merge846(
.A_N(net457),
.B(net472),
.X(net720)
);

sky130_fd_sc_hd__nand2b_2 merge847(
.A_N(net636),
.B(net620),
.Y(net721)
);

sky130_fd_sc_hd__dfsbp_1 merge848(
.D(net648),
.SET_B(net78),
.CLK(clk),
.Q(net723),
.Q_N(net722)
);

sky130_fd_sc_hd__dfsbp_2 merge849(
.D(net652),
.SET_B(net661),
.CLK(clk),
.Q(net725),
.Q_N(net724)
);

sky130_fd_sc_hd__dfstp_1 merge850(
.D(net51),
.SET_B(net676),
.CLK(clk),
.Q(net726)
);

sky130_fd_sc_hd__dfstp_2 merge851(
.D(net242),
.SET_B(net247),
.CLK(clk),
.Q(net727)
);

sky130_fd_sc_hd__dfstp_4 merge852(
.D(net657),
.SET_B(net662),
.CLK(clk),
.Q(net728)
);

sky130_fd_sc_hd__and2_1 merge853(
.A(net502),
.B(net506),
.X(net729)
);

sky130_fd_sc_hd__nor2b_2 merge854(
.A(net328),
.B_N(net344),
.Y(net730)
);

sky130_fd_sc_hd__nor2_1 merge855(
.A(net599),
.B(net603),
.Y(net731)
);

sky130_fd_sc_hd__or2b_4 merge856(
.A(net147),
.B_N(net150),
.X(net732)
);

sky130_fd_sc_hd__nor2b_4 merge857(
.A(net177),
.B_N(net637),
.Y(net733)
);

sky130_fd_sc_hd__dlrbn_1 merge858(
.D(net160),
.RESET_B(net165),
.GATE_N(clk),
.Q(net735),
.Q_N(net734)
);

sky130_fd_sc_hd__dlrbn_2 merge859(
.D(net422),
.RESET_B(net666),
.GATE_N(clk),
.Q(net737),
.Q_N(net736)
);

sky130_fd_sc_hd__nor2_4 merge860(
.A(net289),
.B(net276),
.Y(net738)
);

sky130_fd_sc_hd__nand2_4 merge861(
.A(net362),
.B(net477),
.Y(net739)
);

sky130_fd_sc_hd__nand2_1 merge862(
.A(net364),
.B(net368),
.Y(net740)
);

sky130_fd_sc_hd__nor2b_1 merge863(
.A(net589),
.B_N(net633),
.Y(net741)
);

sky130_fd_sc_hd__and2b_1 merge864(
.A_N(net409),
.B(net401),
.X(net742)
);

sky130_fd_sc_hd__nand2b_1 merge865(
.A_N(net476),
.B(net617),
.Y(net743)
);

sky130_fd_sc_hd__dlrbp_1 merge866(
.D(net298),
.RESET_B(net678),
.GATE(clk),
.Q(out45),
.Q_N(net744)
);

sky130_fd_sc_hd__and2_4 merge867(
.A(net514),
.B(net407),
.X(net745)
);

sky130_fd_sc_hd__dlrbp_2 merge868(
.D(net687),
.RESET_B(net696),
.GATE(clk),
.Q(net747),
.Q_N(net746)
);

sky130_fd_sc_hd__dlrtn_1 merge869(
.D(net167),
.RESET_B(net698),
.GATE_N(clk),
.Q(net748)
);

sky130_fd_sc_hd__dlrtn_2 merge870(
.D(net742),
.RESET_B(net665),
.GATE_N(clk),
.Q(out33)
);

sky130_fd_sc_hd__dlrtn_4 merge871(
.D(net671),
.RESET_B(net102),
.GATE_N(clk),
.Q(net749)
);

sky130_fd_sc_hd__and2_1 merge872(
.A(net592),
.B(net586),
.X(net750)
);

sky130_fd_sc_hd__dlrtp_1 merge873(
.D(net170),
.RESET_B(net658),
.GATE(clk),
.Q(net751)
);

sky130_fd_sc_hd__nor2b_1 merge874(
.A(net604),
.B_N(net616),
.Y(net752)
);

sky130_fd_sc_hd__nor2b_2 merge875(
.A(net625),
.B_N(net508),
.Y(net753)
);

sky130_fd_sc_hd__nor2_4 merge876(
.A(net721),
.B(net521),
.Y(net754)
);

sky130_fd_sc_hd__dlrtp_2 merge877(
.D(net664),
.RESET_B(net667),
.GATE(clk),
.Q(net755)
);

sky130_fd_sc_hd__dlrtp_4 merge878(
.D(net454),
.RESET_B(net741),
.GATE(clk),
.Q(net756)
);

sky130_fd_sc_hd__nor2_1 merge879(
.A(net605),
.B(net520),
.Y(net757)
);

sky130_fd_sc_hd__and2b_1 merge880(
.A_N(net694),
.B(net701),
.X(net758)
);

sky130_fd_sc_hd__edfxbp_1 merge881(
.D(net650),
.DE(net169),
.CLK(clk),
.Q(net760),
.Q_N(net759)
);

sky130_fd_sc_hd__edfxtp_1 merge882(
.D(net451),
.DE(net693),
.CLK(clk),
.Q(net761)
);

sky130_fd_sc_hd__sdlclkp_1 merge883(
.GATE(net677),
.SCE(net699),
.CLK(clk),
.GCLK(net762)
);

sky130_fd_sc_hd__and2b_4 merge884(
.A_N(net518),
.B(net517),
.X(net763)
);

sky130_fd_sc_hd__and2b_4 merge885(
.A_N(net507),
.B(net509),
.X(net764)
);

sky130_fd_sc_hd__nand2b_4 merge886(
.A_N(net606),
.B(net516),
.Y(net765)
);

sky130_fd_sc_hd__sdlclkp_2 merge887(
.GATE(net683),
.SCE(net685),
.CLK(clk),
.GCLK(net766)
);

sky130_fd_sc_hd__sdlclkp_4 merge888(
.GATE(net641),
.SCE(net697),
.CLK(clk),
.GCLK(net767)
);

sky130_fd_sc_hd__dfrbp_1 merge889(
.D(net740),
.RESET_B(net673),
.CLK(clk),
.Q(out35),
.Q_N(net768)
);

sky130_fd_sc_hd__dfrbp_2 merge890(
.D(net220),
.RESET_B(net659),
.CLK(clk),
.Q(net770),
.Q_N(net769)
);

sky130_fd_sc_hd__dfrtn_1 merge891(
.D(net639),
.RESET_B(net692),
.CLK_N(clk),
.Q(net771)
);

sky130_fd_sc_hd__dfrtp_1 merge892(
.D(net287),
.RESET_B(net668),
.CLK(clk),
.Q(net772)
);

sky130_fd_sc_hd__dfrtp_2 merge893(
.D(net675),
.RESET_B(net645),
.CLK(clk),
.Q(net773)
);

sky130_fd_sc_hd__nand2b_1 merge894(
.A_N(net511),
.B(net764),
.Y(net774)
);

sky130_fd_sc_hd__dfrtp_4 merge895(
.D(net79),
.RESET_B(net713),
.CLK(clk),
.Q(net775)
);

sky130_fd_sc_hd__nor2b_4 merge896(
.A(net288),
.B_N(net285),
.Y(net776)
);

sky130_fd_sc_hd__and2_0 merge897(
.A(net609),
.B(net607),
.X(net777)
);

sky130_fd_sc_hd__dfsbp_1 merge898(
.D(net679),
.SET_B(net691),
.CLK(clk),
.Q(net779),
.Q_N(net778)
);

sky130_fd_sc_hd__dfsbp_2 merge899(
.D(net684),
.SET_B(net695),
.CLK(clk),
.Q(net781),
.Q_N(net780)
);

sky130_fd_sc_hd__dfstp_1 merge900(
.D(net688),
.SET_B(net739),
.CLK(clk),
.Q(net782)
);

sky130_fd_sc_hd__dfstp_2 merge901(
.D(net774),
.SET_B(net745),
.CLK(clk),
.Q(net783)
);

sky130_fd_sc_hd__dfstp_4 merge902(
.D(net653),
.SET_B(net753),
.CLK(clk),
.Q(net784)
);

sky130_fd_sc_hd__dlrbn_1 merge903(
.D(net708),
.RESET_B(net496),
.GATE_N(clk),
.Q(net786),
.Q_N(net785)
);

sky130_fd_sc_hd__dlrbn_2 merge904(
.D(net338),
.RESET_B(net356),
.GATE_N(clk),
.Q(net788),
.Q_N(net787)
);

sky130_fd_sc_hd__dlrbp_1 merge905(
.D(net754),
.RESET_B(net410),
.GATE(clk),
.Q(net789),
.Q_N(out24)
);

sky130_fd_sc_hd__dlrbp_2 merge906(
.D(net681),
.RESET_B(net396),
.GATE(clk),
.Q(net790),
.Q_N(out40)
);

sky130_fd_sc_hd__dlrtn_1 merge907(
.D(net743),
.RESET_B(net765),
.GATE_N(clk),
.Q(net791)
);

sky130_fd_sc_hd__dlrtn_2 merge908(
.D(net776),
.RESET_B(net719),
.GATE_N(clk),
.Q(net792)
);

sky130_fd_sc_hd__dlrtn_4 merge909(
.D(net260),
.RESET_B(net709),
.GATE_N(clk),
.Q(net793)
);

sky130_fd_sc_hd__dlrtp_1 merge910(
.D(net394),
.RESET_B(net399),
.GATE(clk),
.Q(out41)
);

sky130_fd_sc_hd__dlrtp_2 merge911(
.D(net321),
.RESET_B(net720),
.GATE(clk),
.Q(net794)
);

sky130_fd_sc_hd__dlrtp_4 merge912(
.D(net717),
.RESET_B(net405),
.GATE(clk),
.Q(out37)
);

sky130_fd_sc_hd__edfxbp_1 merge913(
.D(net646),
.DE(net682),
.CLK(clk),
.Q(net796),
.Q_N(net795)
);

sky130_fd_sc_hd__edfxtp_1 merge914(
.D(net660),
.DE(net750),
.CLK(clk),
.Q(net797)
);

sky130_fd_sc_hd__sdlclkp_1 merge915(
.GATE(net680),
.SCE(net654),
.CLK(clk),
.GCLK(net798)
);

sky130_fd_sc_hd__sdlclkp_2 merge916(
.GATE(net389),
.SCE(net632),
.CLK(clk),
.GCLK(net799)
);

sky130_fd_sc_hd__sdlclkp_4 merge917(
.GATE(net672),
.SCE(net647),
.CLK(clk),
.GCLK(net800)
);

sky130_fd_sc_hd__dfrbp_1 merge918(
.D(net649),
.RESET_B(net757),
.CLK(clk),
.Q(net802),
.Q_N(net801)
);

sky130_fd_sc_hd__dfrbp_2 merge919(
.D(net484),
.RESET_B(net715),
.CLK(clk),
.Q(net804),
.Q_N(net803)
);

sky130_fd_sc_hd__dfrtn_1 merge920(
.D(net642),
.RESET_B(net631),
.CLK_N(clk),
.Q(net805)
);

sky130_fd_sc_hd__dfrtp_1 merge921(
.D(net354),
.RESET_B(net730),
.CLK(clk),
.Q(net806)
);

sky130_fd_sc_hd__dfrtp_2 merge922(
.D(net689),
.RESET_B(net478),
.CLK(clk),
.Q(out2)
);

sky130_fd_sc_hd__dfrtp_4 merge923(
.D(net700),
.RESET_B(net752),
.CLK(clk),
.Q(net807)
);

sky130_fd_sc_hd__dfsbp_1 merge924(
.D(net705),
.SET_B(net763),
.CLK(clk),
.Q(net809),
.Q_N(net808)
);

sky130_fd_sc_hd__dfsbp_2 merge925(
.D(net729),
.SET_B(net515),
.CLK(clk),
.Q(net811),
.Q_N(net810)
);

sky130_fd_sc_hd__dfstp_1 merge926(
.D(net777),
.SET_B(net486),
.CLK(clk),
.Q(net812)
);

sky130_fd_sc_hd__dfstp_2 merge927(
.D(net731),
.SET_B(net690),
.CLK(clk),
.Q(net813)
);

sky130_fd_sc_hd__dfstp_4 merge928(
.D(net738),
.SET_B(net711),
.CLK(clk),
.Q(out48)
);

sky130_fd_sc_hd__dlrbn_1 merge929(
.D(net191),
.RESET_B(net758),
.GATE_N(clk),
.Q(net815),
.Q_N(net814)
);

sky130_fd_sc_hd__dlrbn_2 merge930(
.D(net619),
.RESET_B(net601),
.GATE_N(clk),
.Q(net817),
.Q_N(net816)
);

sky130_fd_sc_hd__dlrbp_1 merge931(
.D(net367),
.RESET_B(net716),
.GATE(clk),
.Q(out43),
.Q_N(net818)
);

sky130_fd_sc_hd__dlrbp_2 merge932(
.D(net732),
.RESET_B(net733),
.GATE(clk),
.Q(net819),
.Q_N(out14)
);

sky130_fd_sc_hd__dfxbp_1 s933(
.D(net24),
.CLK(clk),
.Q(net821),
.Q_N(net820)
);

sky130_fd_sc_hd__dfxbp_2 s934(
.D(net26),
.CLK(clk),
.Q(net823),
.Q_N(net822)
);

sky130_fd_sc_hd__dfxtp_1 s935(
.D(net43),
.CLK(clk),
.Q(net824)
);

sky130_fd_sc_hd__dfxtp_2 s936(
.D(net47),
.CLK(clk),
.Q(net825)
);

sky130_fd_sc_hd__dfxtp_4 s937(
.D(net80),
.CLK(clk),
.Q(net826)
);

sky130_fd_sc_hd__dlclkp_1 s938(
.GATE(net81),
.CLK(clk),
.GCLK(net827)
);

sky130_fd_sc_hd__dlclkp_2 s939(
.GATE(net82),
.CLK(clk),
.GCLK(net828)
);

sky130_fd_sc_hd__dlclkp_4 s940(
.GATE(net83),
.CLK(clk),
.GCLK(net829)
);

sky130_fd_sc_hd__dlxbn_1 s941(
.D(net99),
.GATE_N(clk),
.Q(net831),
.Q_N(net830)
);

sky130_fd_sc_hd__dlxbn_2 s942(
.D(net125),
.GATE_N(clk),
.Q(net833),
.Q_N(net832)
);

sky130_fd_sc_hd__dlxbp_1 s943(
.D(net127),
.GATE(clk),
.Q(net835),
.Q_N(net834)
);

sky130_fd_sc_hd__dlxtn_1 s944(
.D(net166),
.GATE_N(clk),
.Q(net836)
);

sky130_fd_sc_hd__dlxtn_2 s945(
.D(net171),
.GATE_N(clk),
.Q(net837)
);

sky130_fd_sc_hd__dlxtn_4 s946(
.D(net200),
.GATE_N(clk),
.Q(net838)
);

sky130_fd_sc_hd__dlxtp_1 s947(
.D(net202),
.GATE(clk),
.Q(net839)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s948(
.D(net246),
.SLEEP_B(clk),
.Q(net840)
);

sky130_fd_sc_hd__dfxbp_1 s949(
.D(net253),
.CLK(clk),
.Q(net842),
.Q_N(net841)
);

sky130_fd_sc_hd__dfxbp_2 s950(
.D(net269),
.CLK(clk),
.Q(out21),
.Q_N(net843)
);

sky130_fd_sc_hd__dfxtp_1 s951(
.D(net270),
.CLK(clk),
.Q(net844)
);

sky130_fd_sc_hd__dfxtp_2 s952(
.D(net271),
.CLK(clk),
.Q(net845)
);

sky130_fd_sc_hd__dfxtp_4 s953(
.D(net273),
.CLK(clk),
.Q(net846)
);

sky130_fd_sc_hd__dlclkp_1 s954(
.GATE(net286),
.CLK(clk),
.GCLK(net847)
);

sky130_fd_sc_hd__dlclkp_2 s955(
.GATE(net343),
.CLK(clk),
.GCLK(net848)
);

sky130_fd_sc_hd__dlclkp_4 s956(
.GATE(net346),
.CLK(clk),
.GCLK(net849)
);

sky130_fd_sc_hd__dlxbn_1 s957(
.D(net365),
.GATE_N(clk),
.Q(net851),
.Q_N(net850)
);

sky130_fd_sc_hd__dlxbn_2 s958(
.D(net411),
.GATE_N(clk),
.Q(net853),
.Q_N(net852)
);

sky130_fd_sc_hd__dlxbp_1 s959(
.D(net429),
.GATE(clk),
.Q(net855),
.Q_N(net854)
);

sky130_fd_sc_hd__dlxtn_1 s960(
.D(net431),
.GATE_N(clk),
.Q(net856)
);

sky130_fd_sc_hd__dlxtn_2 s961(
.D(net433),
.GATE_N(clk),
.Q(net857)
);

sky130_fd_sc_hd__dlxtn_4 s962(
.D(net446),
.GATE_N(clk),
.Q(net858)
);

sky130_fd_sc_hd__dlxtp_1 s963(
.D(net449),
.GATE(clk),
.Q(net859)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s964(
.D(net456),
.SLEEP_B(clk),
.Q(net860)
);

sky130_fd_sc_hd__dfxbp_1 s965(
.D(net483),
.CLK(clk),
.Q(net862),
.Q_N(net861)
);

sky130_fd_sc_hd__dfxbp_2 s966(
.D(net487),
.CLK(clk),
.Q(net864),
.Q_N(net863)
);

sky130_fd_sc_hd__dfxtp_1 s967(
.D(net497),
.CLK(clk),
.Q(out10)
);

sky130_fd_sc_hd__dfxtp_2 s968(
.D(net499),
.CLK(clk),
.Q(net865)
);

sky130_fd_sc_hd__dfxtp_4 s969(
.D(net500),
.CLK(clk),
.Q(net866)
);

sky130_fd_sc_hd__dlclkp_1 s970(
.GATE(net503),
.CLK(clk),
.GCLK(net867)
);

sky130_fd_sc_hd__dlclkp_2 s971(
.GATE(net510),
.CLK(clk),
.GCLK(out20)
);

sky130_fd_sc_hd__dlclkp_4 s972(
.GATE(net512),
.CLK(clk),
.GCLK(net868)
);

sky130_fd_sc_hd__dlxbn_1 s973(
.D(net522),
.GATE_N(clk),
.Q(net870),
.Q_N(net869)
);

sky130_fd_sc_hd__dlxbn_2 s974(
.D(net535),
.GATE_N(clk),
.Q(net872),
.Q_N(net871)
);

sky130_fd_sc_hd__dlxbp_1 s975(
.D(net563),
.GATE(clk),
.Q(net874),
.Q_N(net873)
);

sky130_fd_sc_hd__dlxtn_1 s976(
.D(net568),
.GATE_N(clk),
.Q(net875)
);

sky130_fd_sc_hd__dlxtn_2 s977(
.D(net569),
.GATE_N(clk),
.Q(net876)
);

sky130_fd_sc_hd__dlxtn_4 s978(
.D(net579),
.GATE_N(clk),
.Q(net877)
);

sky130_fd_sc_hd__dlxtp_1 s979(
.D(net588),
.GATE(clk),
.Q(net878)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s980(
.D(net590),
.SLEEP_B(clk),
.Q(net879)
);

sky130_fd_sc_hd__dfxbp_1 s981(
.D(net594),
.CLK(clk),
.Q(net881),
.Q_N(net880)
);

sky130_fd_sc_hd__dfxbp_2 s982(
.D(net595),
.CLK(clk),
.Q(net883),
.Q_N(net882)
);

sky130_fd_sc_hd__dfxtp_1 s983(
.D(net602),
.CLK(clk),
.Q(net884)
);

sky130_fd_sc_hd__dfxtp_2 s984(
.D(net608),
.CLK(clk),
.Q(net885)
);

sky130_fd_sc_hd__dfxtp_4 s985(
.D(net610),
.CLK(clk),
.Q(net886)
);

sky130_fd_sc_hd__dlclkp_1 s986(
.GATE(net611),
.CLK(clk),
.GCLK(net887)
);

sky130_fd_sc_hd__dlclkp_2 s987(
.GATE(net612),
.CLK(clk),
.GCLK(net888)
);

sky130_fd_sc_hd__dlclkp_4 s988(
.GATE(net615),
.CLK(clk),
.GCLK(net889)
);

sky130_fd_sc_hd__dlxbn_1 s989(
.D(net621),
.GATE_N(clk),
.Q(net891),
.Q_N(net890)
);

sky130_fd_sc_hd__dlxbn_2 s990(
.D(net627),
.GATE_N(clk),
.Q(net893),
.Q_N(net892)
);

sky130_fd_sc_hd__dlxbp_1 s991(
.D(net629),
.GATE(clk),
.Q(net895),
.Q_N(net894)
);

sky130_fd_sc_hd__dlxtn_1 s992(
.D(net686),
.GATE_N(clk),
.Q(net896)
);

sky130_fd_sc_hd__dlxtn_2 s993(
.D(net702),
.GATE_N(clk),
.Q(net897)
);


endmodule
