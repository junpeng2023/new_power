module netlist_0 (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input in26,
	input in27,
	input in28,
	input in29,
	input in30,
	input in31,
	input in32,
	input in33,
	input in34,
	input in35,
	input in36,
	input in37,
	input in38,
	input in39,
	input in40,
	input in41,
	input in42,
	input in43,
	input in44,
	input in45,
	input in46,
	input in47,
	input in48,
	input in49,
	input in50,
	input in51,
	input in52,
	input in53,
	input in54,
	input in55,
	input in56,
	input in57,
	input in58,
	input in59,
	input in60,
	input in61,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25,
	output out26,
	output out27,
	output out28,
	output out29,
	output out30,
	output out31,
	output out32,
	output out33,
	output out34,
	output out35,
	output out36,
	output out37,
	output out38,
	output out39,
	output out40,
	output out41,
	output out42,
	output out43,
	output out44,
	output out45,
	output out46,
	output out47,
	output out48,
	output out49,
	output out50,
	output out51,
	output out52,
	output out53,
	output out54,
	output out55,
	output out56,
	output out57,
	output out58,
	output out59,
	output out60,
	output out61
);


wire clk;
wire net695;
wire net694;
wire net693;
wire net692;
wire net690;
wire net687;
wire net686;
wire net685;
wire net684;
wire net683;
wire net680;
wire net678;
wire net676;
wire net671;
wire net669;
wire net668;
wire net370;
wire net667;
wire net664;
wire net659;
wire out54;
wire in6;
wire net656;
wire net652;
wire net622;
wire net651;
wire net304;
wire net645;
wire net641;
wire net637;
wire net632;
wire net665;
wire net631;
wire net629;
wire net74;
wire net628;
wire net3;
wire net627;
wire net447;
wire net626;
wire net624;
wire net506;
wire net623;
wire net620;
wire in49;
wire net619;
wire net46;
wire net615;
wire net100;
wire net347;
wire net288;
wire net614;
wire net165;
wire net613;
wire net20;
wire net612;
wire net638;
wire net428;
wire net610;
wire out25;
wire net608;
wire net1;
wire net424;
wire net606;
wire net605;
wire net604;
wire net603;
wire net602;
wire net596;
wire out52;
wire net384;
wire net482;
wire net595;
wire net592;
wire net588;
wire net587;
wire in4;
wire net583;
wire net582;
wire net158;
wire net584;
wire net581;
wire net336;
wire net579;
wire net577;
wire net576;
wire net209;
wire net569;
wire in41;
wire net567;
wire in30;
wire net566;
wire net565;
wire net39;
wire net562;
wire net559;
wire net556;
wire net647;
wire net555;
wire net159;
wire net635;
wire net554;
wire net553;
wire net552;
wire net551;
wire in55;
wire net550;
wire net544;
wire net539;
wire net534;
wire net532;
wire net271;
wire net530;
wire net617;
wire net306;
wire net537;
wire net369;
wire net528;
wire net525;
wire net523;
wire net520;
wire net519;
wire net516;
wire net672;
wire net514;
wire net18;
wire out34;
wire net512;
wire net78;
wire net508;
wire net504;
wire net679;
wire out57;
wire net503;
wire net224;
wire net573;
wire net499;
wire net674;
wire net496;
wire out17;
wire net495;
wire net494;
wire net179;
wire in39;
wire net453;
wire net493;
wire net472;
wire net492;
wire net479;
wire net491;
wire net295;
wire net490;
wire net489;
wire net487;
wire net486;
wire net478;
wire out20;
wire net474;
wire net473;
wire out13;
wire net468;
wire net540;
wire net202;
wire net465;
wire out7;
wire net462;
wire net469;
wire net471;
wire net461;
wire net546;
wire net460;
wire net454;
wire net648;
wire net452;
wire net449;
wire net448;
wire net498;
wire net446;
wire net691;
wire net88;
wire net444;
wire in59;
wire net110;
wire net442;
wire out15;
wire net441;
wire net609;
wire net440;
wire net128;
wire net439;
wire net147;
wire out21;
wire net438;
wire net433;
wire net432;
wire net419;
wire net431;
wire net430;
wire net618;
wire net429;
wire net427;
wire net426;
wire net673;
wire net425;
wire net423;
wire net183;
wire net531;
wire net421;
wire net52;
wire net170;
wire net420;
wire net450;
wire net418;
wire net415;
wire net414;
wire net276;
wire net413;
wire net252;
wire net330;
wire net412;
wire net411;
wire net410;
wire net409;
wire net407;
wire out19;
wire net406;
wire net662;
wire net405;
wire net607;
wire net526;
wire net404;
wire net29;
wire net403;
wire net383;
wire net663;
wire net402;
wire net106;
wire net572;
wire net401;
wire net399;
wire net398;
wire net476;
wire net396;
wire net391;
wire net443;
wire net557;
wire net345;
wire net527;
wire net488;
wire net390;
wire net475;
wire net408;
wire out26;
wire out5;
wire net646;
wire net389;
wire net513;
wire net501;
wire out14;
wire net388;
wire net545;
wire net387;
wire net634;
wire net386;
wire net385;
wire net184;
wire net131;
wire net380;
wire net379;
wire net260;
wire net616;
wire net378;
wire out37;
wire net543;
wire net38;
wire net377;
wire net376;
wire net625;
wire net373;
wire net598;
wire net374;
wire net372;
wire net371;
wire net368;
wire net416;
wire net41;
wire net104;
wire net8;
wire out33;
wire net367;
wire net366;
wire net365;
wire net364;
wire net363;
wire net360;
wire net397;
wire net357;
wire net356;
wire net510;
wire net355;
wire net590;
wire net507;
wire net351;
wire net350;
wire net547;
wire net511;
wire net451;
wire net13;
wire net343;
wire net89;
wire net666;
wire net340;
wire net339;
wire net337;
wire net458;
wire net538;
wire net244;
wire net334;
wire net333;
wire net332;
wire net331;
wire out32;
wire net677;
wire net517;
wire net328;
wire net327;
wire net119;
wire net325;
wire net324;
wire net321;
wire net535;
wire net320;
wire net542;
wire net139;
wire net318;
wire out9;
wire net335;
wire net315;
wire net313;
wire net505;
wire net199;
wire out27;
wire net294;
wire net319;
wire net312;
wire net309;
wire net308;
wire net352;
wire net307;
wire net305;
wire net291;
wire net303;
wire net301;
wire net298;
wire net459;
wire net463;
wire net0;
wire net297;
wire net296;
wire in24;
wire net358;
wire net127;
wire net293;
wire net594;
wire out39;
wire net292;
wire net500;
wire net445;
wire net230;
wire out22;
wire net201;
wire net422;
wire net289;
wire in25;
wire out58;
wire net589;
wire net278;
wire out49;
wire net274;
wire net643;
wire net273;
wire net142;
wire out10;
wire net272;
wire net114;
wire net270;
wire in17;
wire net267;
wire in8;
wire net30;
wire out36;
wire net644;
wire net266;
wire out6;
wire net521;
wire net353;
wire net280;
wire net102;
wire net151;
wire net275;
wire net264;
wire net657;
wire net591;
wire net196;
wire net262;
wire net217;
wire net261;
wire net21;
wire net257;
wire net689;
wire net44;
wire net117;
wire net62;
wire net109;
wire net254;
wire net203;
wire net253;
wire net188;
wire net207;
wire out16;
wire net249;
wire net66;
wire net247;
wire net245;
wire net10;
wire in40;
wire net243;
wire in26;
wire net661;
wire net194;
wire net241;
wire in29;
wire net240;
wire out42;
wire net238;
wire net234;
wire net232;
wire out12;
wire net226;
wire net568;
wire net375;
wire net223;
wire net524;
wire net575;
wire net382;
wire net548;
wire net259;
wire net222;
wire net31;
wire net219;
wire net578;
wire net210;
wire net326;
wire net213;
wire net208;
wire net649;
wire net205;
wire net633;
wire net122;
wire net197;
wire net483;
wire net193;
wire net192;
wire net190;
wire net630;
wire in20;
wire net189;
wire net246;
wire net186;
wire net152;
wire net126;
wire net113;
wire net284;
wire net655;
wire net563;
wire net464;
wire net549;
wire net182;
wire net310;
wire net180;
wire net342;
wire net17;
wire net437;
wire out44;
wire net580;
wire net133;
wire net175;
wire net80;
wire net173;
wire net195;
wire net395;
wire net172;
wire in37;
wire net518;
wire net381;
wire net218;
wire net300;
wire net169;
wire net485;
wire net344;
wire net168;
wire net111;
wire net124;
wire net242;
wire net290;
wire net227;
wire out47;
wire net153;
wire net286;
wire net167;
wire net509;
wire net58;
wire net221;
wire net166;
wire net269;
wire out3;
wire net97;
wire net434;
wire net204;
wire net200;
wire net621;
wire net162;
wire out60;
wire net497;
wire out45;
wire net161;
wire net285;
wire net160;
wire net636;
wire net311;
wire net417;
wire net302;
wire out8;
wire net150;
wire net149;
wire net148;
wire net178;
wire net239;
wire net144;
wire net322;
wire net688;
wire net299;
wire net143;
wire net141;
wire net140;
wire net283;
wire net83;
wire net287;
wire net561;
wire out29;
wire net137;
wire net136;
wire net456;
wire net135;
wire net255;
wire net157;
wire net177;
wire net349;
wire out51;
wire net134;
wire net250;
wire net225;
wire net132;
wire net130;
wire net642;
wire net268;
wire in7;
wire net400;
wire net82;
wire net2;
wire net123;
wire out18;
wire net481;
wire net120;
wire net392;
wire out0;
wire net164;
wire net282;
wire net71;
wire net229;
wire in43;
wire net108;
wire net107;
wire in12;
wire net103;
wire net6;
wire net457;
wire out50;
wire net348;
wire net341;
wire in52;
wire net96;
wire net466;
wire net118;
wire net94;
wire net90;
wire net174;
wire net277;
wire net639;
wire net81;
wire in10;
wire net156;
wire net361;
wire net115;
wire net670;
wire in18;
wire net27;
wire net34;
wire net258;
wire out40;
wire net585;
wire net79;
wire net231;
wire net329;
wire net212;
wire net653;
wire in5;
wire net14;
wire net77;
wire net600;
wire net236;
wire net76;
wire in42;
wire net354;
wire in38;
wire net198;
wire net467;
wire net101;
wire net9;
wire net75;
wire net571;
wire net73;
wire net60;
wire net564;
wire net154;
wire net84;
wire in46;
wire net85;
wire net72;
wire net116;
wire net69;
wire net98;
wire net522;
wire net436;
wire net541;
wire net323;
wire net15;
wire net279;
wire net64;
wire net63;
wire net681;
wire net61;
wire net682;
wire net237;
wire net59;
wire net228;
wire net675;
wire net56;
wire out53;
wire net55;
wire net640;
wire net50;
wire net67;
wire net92;
wire net25;
wire net214;
wire net53;
wire in48;
wire in31;
wire net129;
wire net65;
wire net660;
wire net359;
wire out28;
wire net597;
wire out55;
wire net185;
wire net155;
wire net338;
wire net599;
wire net112;
wire net650;
wire net560;
wire net45;
wire net502;
wire net235;
wire net49;
wire in50;
wire net215;
wire net484;
wire net346;
wire net4;
wire net43;
wire net99;
wire net211;
wire net145;
wire net574;
wire net26;
wire net23;
wire out1;
wire net233;
wire net33;
wire net187;
wire in13;
wire net586;
wire net533;
wire net32;
wire net125;
wire net19;
wire in15;
wire net163;
wire in19;
wire net70;
wire net48;
wire net28;
wire net570;
wire out2;
wire in0;
wire net24;
wire out59;
wire net176;
wire out23;
wire net470;
wire in33;
wire net40;
wire in60;
wire net435;
wire net16;
wire net558;
wire in1;
wire net265;
wire net22;
wire net263;
wire net5;
wire net206;
wire in58;
wire in61;
wire in56;
wire net171;
wire in23;
wire out4;
wire net42;
wire net91;
wire in57;
wire net281;
wire net54;
wire in54;
wire out43;
wire in53;
wire out11;
wire net138;
wire out24;
wire in35;
wire in34;
wire net593;
wire in45;
wire net393;
wire net256;
wire net87;
wire net181;
wire net7;
wire net216;
wire net455;
wire in28;
wire in44;
wire net601;
wire out35;
wire in32;
wire net47;
wire net12;
wire in27;
wire net536;
wire net37;
wire in9;
wire net654;
wire net611;
wire net515;
wire net362;
wire in16;
wire net191;
wire out46;
wire net35;
wire net220;
wire in22;
wire net68;
wire in14;
wire net529;
wire in21;
wire net248;
wire net477;
wire out38;
wire out56;
wire net57;
wire net480;
wire net86;
wire net317;
wire in51;
wire net93;
wire in47;
wire in2;
wire net658;
wire net105;
wire in11;
wire net51;
wire out30;
wire in36;
wire net316;
wire out31;
wire net36;
wire net95;
wire net121;
wire net146;
wire net251;
wire net11;
wire net394;
wire net314;
wire in3;
sky130_fd_sc_hd__o2111ai_1 c62(
.A1(in61),
.A2(in40),
.B1(in29),
.C1(in50),
.D1(in27),
.Y(net0)
);

sky130_fd_sc_hd__mux4_1 c63(
.A0(net0),
.A1(in44),
.A2(in47),
.A3(net2),
.S0(in60),
.S1(in50),
.X(out0)
);

sky130_fd_sc_hd__mux4_1 c64(
.A0(in34),
.A1(in47),
.A2(in27),
.A3(in44),
.S0(in52),
.S1(net0),
.X(net1)
);

sky130_fd_sc_hd__nand3b_4 c65(
.A_N(in26),
.B(in19),
.C(in34),
.Y(net2)
);

sky130_fd_sc_hd__nor2b_4 c66(
.A(in47),
.B_N(in59),
.Y(net3)
);

sky130_fd_sc_hd__or2b_1 c67(
.A(in55),
.B_N(in0),
.X(net4)
);

sky130_fd_sc_hd__or2b_2 c68(
.A(in27),
.B_N(net3),
.X(net5)
);

sky130_fd_sc_hd__nand2_2 c69(
.A(in39),
.B(net4),
.Y(net6)
);

sky130_fd_sc_hd__nand2b_4 c70(
.A_N(in50),
.B(net4),
.Y(net7)
);

sky130_fd_sc_hd__nand2b_4 c71(
.A_N(in57),
.B(in52),
.Y(net8)
);

sky130_fd_sc_hd__nand2b_2 c72(
.A_N(net6),
.B(net8),
.Y(net9)
);

sky130_fd_sc_hd__nand2_4 c73(
.A(net1),
.B(net7),
.Y(net10)
);

sky130_fd_sc_hd__nand2_1 c74(
.A(net9),
.B(net10),
.Y(net11)
);

sky130_fd_sc_hd__or2b_2 c75(
.A(in44),
.B_N(net4),
.X(net12)
);

sky130_fd_sc_hd__and2b_2 c76(
.A_N(net7),
.B(net9),
.X(net13)
);

sky130_fd_sc_hd__nand3b_1 c77(
.A_N(in19),
.B(in50),
.C(net7),
.Y(net14)
);

sky130_fd_sc_hd__nand2_1 c78(
.A(net11),
.B(net12),
.Y(net15)
);

sky130_fd_sc_hd__nor2_4 c79(
.A(in52),
.B(net15),
.Y(out56)
);

sky130_fd_sc_hd__or2_1 c80(
.A(net15),
.B(net14),
.X(net16)
);

sky130_fd_sc_hd__or2b_1 c81(
.A(net12),
.B_N(in45),
.X(net17)
);

sky130_fd_sc_hd__nor2b_1 c82(
.A(net16),
.B_N(net8),
.Y(net18)
);

sky130_fd_sc_hd__and2b_2 c83(
.A_N(in45),
.B(net3),
.X(net19)
);

sky130_fd_sc_hd__nor2b_1 c84(
.A(net19),
.B_N(net17),
.Y(net20)
);

sky130_fd_sc_hd__or2_1 c85(
.A(net13),
.B(net20),
.X(net21)
);

sky130_fd_sc_hd__or3_2 c86(
.A(net17),
.B(net16),
.C(net14),
.X(net22)
);

sky130_fd_sc_hd__nor2b_1 c87(
.A(net5),
.B_N(net22),
.Y(net23)
);

sky130_fd_sc_hd__or2b_2 c88(
.A(in28),
.B_N(net22),
.X(net24)
);

sky130_fd_sc_hd__or2b_4 c89(
.A(in29),
.B_N(in49),
.X(net25)
);

sky130_fd_sc_hd__nand2b_4 c90(
.A_N(net24),
.B(net14),
.Y(net26)
);

sky130_fd_sc_hd__nand3_2 c91(
.A(in61),
.B(net2),
.C(in28),
.Y(net27)
);

sky130_fd_sc_hd__nor2b_4 c92(
.A(net26),
.B_N(net24),
.Y(net28)
);

sky130_fd_sc_hd__nand2_2 c93(
.A(net28),
.B(net22),
.Y(net29)
);

sky130_fd_sc_hd__or2_1 c94(
.A(net27),
.B(net24),
.X(net30)
);

sky130_fd_sc_hd__nor2_2 c95(
.A(in49),
.B(net28),
.Y(net31)
);

sky130_fd_sc_hd__nor2_4 c96(
.A(net31),
.B(net28),
.Y(net32)
);

sky130_fd_sc_hd__and2b_2 c97(
.A_N(net26),
.B(net32),
.X(net33)
);

sky130_fd_sc_hd__nand2b_1 c98(
.A_N(net33),
.B(net26),
.Y(net34)
);

sky130_fd_sc_hd__and2b_4 c99(
.A_N(net32),
.B(net34),
.X(out1)
);

sky130_fd_sc_hd__or2_1 c100(
.A(net30),
.B(net31),
.X(net35)
);

sky130_fd_sc_hd__and2b_1 c101(
.A_N(net28),
.B(net26),
.X(net36)
);

sky130_fd_sc_hd__nand2_2 c102(
.A(in20),
.B(net13),
.Y(net37)
);

sky130_fd_sc_hd__or2b_2 c103(
.A(in31),
.B_N(net34),
.X(net38)
);

sky130_fd_sc_hd__nand2_2 c104(
.A(net3),
.B(net32),
.Y(net39)
);

sky130_fd_sc_hd__inv_1 c105(
.Y(net40)
);

sky130_fd_sc_hd__or3_2 c106(
.A(net37),
.B(net26),
.C(net34),
.X(net41)
);

sky130_fd_sc_hd__dlygate4sd1_1 c107(
.A(net619),
.X(net42)
);

sky130_fd_sc_hd__or3_4 c108(
.A(net37),
.B(net36),
.C(net42),
.X(net43)
);

sky130_fd_sc_hd__nor2_1 c109(
.A(net36),
.B(net42),
.Y(net44)
);

sky130_fd_sc_hd__inv_16 c110(
.A(net636),
.Y(net45)
);

sky130_fd_sc_hd__nor2_2 c111(
.A(in0),
.B(net13),
.Y(net46)
);

sky130_fd_sc_hd__nand2_4 c112(
.A(net13),
.B(net45),
.Y(out27)
);

sky130_fd_sc_hd__and2b_1 c113(
.A_N(net14),
.B(net43),
.X(out28)
);

sky130_fd_sc_hd__or2_2 c114(
.A(in48),
.B(in38),
.X(out31)
);

sky130_fd_sc_hd__nand2b_2 c115(
.A_N(net35),
.B(out56),
.Y(out23)
);

sky130_fd_sc_hd__buf_6 c116(
.A(net635),
.X(net47)
);

sky130_fd_sc_hd__nand2b_1 c117(
.A_N(net45),
.B(net14),
.Y(net48)
);

sky130_fd_sc_hd__buf_8 c118(
.A(net640),
.X(net49)
);

sky130_fd_sc_hd__or2_2 c119(
.A(out0),
.B(net49),
.X(out53)
);

sky130_fd_sc_hd__nor2b_2 c120(
.A(net27),
.B_N(net49),
.Y(net50)
);

sky130_fd_sc_hd__or3b_2 c121(
.A(net47),
.B(net46),
.C_N(net49),
.X(net51)
);

sky130_fd_sc_hd__nor2b_4 c122(
.A(net50),
.B_N(net49),
.Y(net52)
);

sky130_fd_sc_hd__nor3_2 c123(
.A(net48),
.B(net50),
.C(net52),
.Y(net53)
);

sky130_fd_sc_hd__or2b_4 c124(
.A(net51),
.B_N(net49),
.X(out39)
);

sky130_fd_sc_hd__nor2_1 c125(
.A(in48),
.B(out39),
.Y(out40)
);

sky130_fd_sc_hd__nand2_4 c126(
.A(net53),
.B(net46),
.Y(out12)
);

sky130_fd_sc_hd__nor2_2 c127(
.A(net49),
.B(out12),
.Y(net54)
);

sky130_fd_sc_hd__and2b_4 c128(
.A_N(net54),
.B(out40),
.X(net55)
);

sky130_fd_sc_hd__nand3b_4 c129(
.A_N(net46),
.B(net55),
.C(net50),
.Y(net56)
);

sky130_fd_sc_hd__or2b_4 c130(
.A(net54),
.B_N(out39),
.X(net57)
);

sky130_fd_sc_hd__or4bb_4 c131(
.A(net52),
.B(net57),
.C_N(out39),
.D_N(net50),
.X(net58)
);

sky130_fd_sc_hd__or2_1 c132(
.A(in12),
.B(in0),
.X(net59)
);

sky130_fd_sc_hd__nor2b_2 c133(
.A(in2),
.B_N(net59),
.Y(net60)
);

sky130_fd_sc_hd__or2b_2 c134(
.A(in16),
.B_N(net60),
.X(net61)
);

sky130_fd_sc_hd__or2_2 c135(
.A(in21),
.B(in16),
.X(net62)
);

sky130_fd_sc_hd__or3b_4 c136(
.A(in9),
.B(in1),
.C_N(in21),
.X(net63)
);

sky130_fd_sc_hd__and2_4 c137(
.A(net63),
.B(in2),
.X(net64)
);

sky130_fd_sc_hd__or2_4 c138(
.A(in16),
.B(net64),
.X(net65)
);

sky130_fd_sc_hd__nor2_2 c139(
.A(in2),
.B(net65),
.Y(net66)
);

sky130_fd_sc_hd__nand2_1 c140(
.A(net66),
.B(net62),
.Y(net67)
);

sky130_fd_sc_hd__and2_2 c141(
.A(net66),
.B(net67),
.X(net68)
);

sky130_fd_sc_hd__nor2_1 c142(
.A(net67),
.B(net61),
.Y(out22)
);

sky130_fd_sc_hd__and2_0 c143(
.A(net62),
.B(net64),
.X(net69)
);

sky130_fd_sc_hd__nor2b_4 c144(
.A(in11),
.B_N(in8),
.Y(net70)
);

sky130_fd_sc_hd__or2b_1 c145(
.A(net69),
.B_N(net61),
.X(net71)
);

sky130_fd_sc_hd__and2_2 c146(
.A(net68),
.B(net69),
.X(net72)
);

sky130_fd_sc_hd__or4bb_4 c147(
.A(net60),
.B(net62),
.C_N(in18),
.D_N(net59),
.X(net73)
);

sky130_fd_sc_hd__nand2_2 c148(
.A(net62),
.B(net71),
.Y(net74)
);

sky130_fd_sc_hd__or3b_1 c149(
.A(net74),
.B(net64),
.C_N(net69),
.X(net75)
);

sky130_fd_sc_hd__and2b_2 c150(
.A_N(net70),
.B(net71),
.X(net76)
);

sky130_fd_sc_hd__nor2_4 c151(
.A(net76),
.B(net75),
.Y(net77)
);

sky130_fd_sc_hd__o2111a_1 c152(
.A1(net72),
.A2(net73),
.B1(net77),
.C1(net69),
.D1(net59),
.X(net78)
);

sky130_fd_sc_hd__or3_2 c153(
.A(net75),
.B(net78),
.C(net76),
.X(net79)
);

sky130_fd_sc_hd__and2b_4 c154(
.A_N(in32),
.B(in22),
.X(net80)
);

sky130_fd_sc_hd__nand2b_4 c155(
.A_N(in42),
.B(net72),
.Y(net81)
);

sky130_fd_sc_hd__nand2b_4 c156(
.A_N(net61),
.B(net72),
.Y(net82)
);

sky130_fd_sc_hd__nand2b_1 c157(
.A_N(net65),
.B(net72),
.Y(net83)
);

sky130_fd_sc_hd__nor2_2 c158(
.A(in18),
.B(net61),
.Y(net84)
);

sky130_fd_sc_hd__and2b_4 c159(
.A_N(net68),
.B(net80),
.X(net85)
);

sky130_fd_sc_hd__nor2b_4 c160(
.A(in38),
.B_N(out22),
.Y(net86)
);

sky130_fd_sc_hd__and2_0 c161(
.A(net83),
.B(in33),
.X(net87)
);

sky130_fd_sc_hd__nand3_4 c162(
.A(in36),
.B(in31),
.C(net85),
.Y(net88)
);

sky130_fd_sc_hd__or2_2 c163(
.A(net85),
.B(net88),
.X(net89)
);

sky130_fd_sc_hd__or2b_1 c164(
.A(net81),
.B_N(net82),
.X(net90)
);

sky130_fd_sc_hd__or2b_2 c165(
.A(in25),
.B_N(in13),
.X(net91)
);

sky130_fd_sc_hd__nor2b_1 c166(
.A(net86),
.B_N(in41),
.Y(net92)
);

sky130_fd_sc_hd__nand2b_4 c167(
.A_N(net90),
.B(net86),
.Y(net93)
);

sky130_fd_sc_hd__and2_0 c168(
.A(net91),
.B(net87),
.X(net94)
);

sky130_fd_sc_hd__nor3_1 c169(
.A(net82),
.B(net91),
.C(net93),
.Y(net95)
);

sky130_fd_sc_hd__or3b_1 c170(
.A(net95),
.B(in13),
.C_N(net90),
.X(net96)
);

sky130_fd_sc_hd__and3_1 c171(
.A(net94),
.B(net93),
.C(net88),
.X(net97)
);

sky130_fd_sc_hd__and2_1 c172(
.A(net87),
.B(net94),
.X(net98)
);

sky130_fd_sc_hd__or4bb_4 c173(
.A(net98),
.B(net97),
.C_N(net93),
.D_N(net85),
.X(net99)
);

sky130_fd_sc_hd__or3b_1 c174(
.A(net92),
.B(net99),
.C_N(in43),
.X(net100)
);

sky130_fd_sc_hd__mux4_1 c175(
.A0(in41),
.A1(net89),
.A2(net100),
.A3(net98),
.S0(net88),
.S1(net85),
.X(net101)
);

sky130_fd_sc_hd__nand2_4 c176(
.A(net84),
.B(in51),
.Y(net102)
);

sky130_fd_sc_hd__or3b_2 c177(
.A(in13),
.B(net84),
.C_N(net85),
.X(net103)
);

sky130_fd_sc_hd__nand3_1 c178(
.A(in56),
.B(net81),
.C(net103),
.Y(net104)
);

sky130_fd_sc_hd__and2b_4 c179(
.A_N(in46),
.B(net2),
.X(net105)
);

sky130_fd_sc_hd__and3_4 c180(
.A(in37),
.B(in3),
.C(net97),
.X(net106)
);

sky130_fd_sc_hd__mux4_1 c181(
.A0(net103),
.A1(net93),
.A2(in22),
.A3(net78),
.S0(net59),
.S1(in59),
.X(net107)
);

sky130_fd_sc_hd__or2_2 c182(
.A(in30),
.B(net59),
.X(net108)
);

sky130_fd_sc_hd__nand2_4 c183(
.A(net78),
.B(net104),
.Y(net109)
);

sky130_fd_sc_hd__nand2_1 c184(
.A(net108),
.B(net80),
.Y(net110)
);

sky130_fd_sc_hd__and2b_1 c185(
.A_N(in51),
.B(net95),
.X(net111)
);

sky130_fd_sc_hd__nor2_2 c186(
.A(net111),
.B(net106),
.Y(net112)
);

sky130_fd_sc_hd__nor2_2 c187(
.A(in24),
.B(net0),
.Y(net113)
);

sky130_fd_sc_hd__and3b_1 c188(
.A_N(net112),
.B(in51),
.C(net111),
.X(net114)
);

sky130_fd_sc_hd__nor2_2 c189(
.A(net106),
.B(net111),
.Y(net115)
);

sky130_fd_sc_hd__nand2_4 c190(
.A(in3),
.B(in32),
.Y(net116)
);

sky130_fd_sc_hd__or3_2 c191(
.A(net104),
.B(net107),
.C(net110),
.X(net117)
);

sky130_fd_sc_hd__or4bb_4 c192(
.A(in54),
.B(net0),
.C_N(in22),
.D_N(net108),
.X(net118)
);

sky130_fd_sc_hd__or4bb_2 c193(
.A(net115),
.B(net117),
.C_N(net114),
.D_N(net73),
.X(net119)
);

sky130_fd_sc_hd__and2_0 c194(
.A(in40),
.B(net107),
.X(net120)
);

sky130_fd_sc_hd__or3b_2 c195(
.A(net117),
.B(net99),
.C_N(net73),
.X(net121)
);

sky130_fd_sc_hd__or4bb_2 c196(
.A(in60),
.B(net120),
.C_N(net115),
.D_N(net121),
.X(net122)
);

sky130_fd_sc_hd__and3b_2 c197(
.A_N(net120),
.B(in30),
.C(net121),
.X(net123)
);

sky130_fd_sc_hd__or2b_1 c198(
.A(net109),
.B_N(in5),
.X(out46)
);

sky130_fd_sc_hd__and2_0 c199(
.A(net120),
.B(net103),
.X(net124)
);

sky130_fd_sc_hd__or4bb_4 c200(
.A(out46),
.B(net113),
.C_N(net123),
.D_N(net18),
.X(net125)
);

sky130_fd_sc_hd__or3b_1 c201(
.A(in31),
.B(net114),
.C_N(out46),
.X(net126)
);

sky130_fd_sc_hd__nand2_1 c202(
.A(net103),
.B(net85),
.Y(net127)
);

sky130_fd_sc_hd__and2b_4 c203(
.A_N(in22),
.B(net23),
.X(net128)
);

sky130_fd_sc_hd__or3_1 c204(
.A(net127),
.B(out56),
.C(net10),
.X(net129)
);

sky130_fd_sc_hd__nor3b_1 c205(
.A(net12),
.B(net129),
.C_N(net15),
.Y(net130)
);

sky130_fd_sc_hd__clkbuf_2 c206(
.A(net618),
.X(net131)
);

sky130_fd_sc_hd__clkbuf_2 c207(
.A(net618),
.X(out11)
);

sky130_fd_sc_hd__nand2b_4 c208(
.A_N(in8),
.B(out11),
.Y(net132)
);

sky130_fd_sc_hd__nand2_1 c209(
.A(net81),
.B(net129),
.Y(net133)
);

sky130_fd_sc_hd__or3_4 c210(
.A(net73),
.B(net12),
.C(out11),
.X(out43)
);

sky130_fd_sc_hd__inv_16 c211(
.A(net639),
.Y(net134)
);

sky130_fd_sc_hd__or3b_1 c212(
.A(net10),
.B(net129),
.C_N(net103),
.X(net135)
);

sky130_fd_sc_hd__nand2_1 c213(
.A(net133),
.B(out46),
.Y(net136)
);

sky130_fd_sc_hd__sdfrbp_1 c214(
.D(net129),
.RESET_B(net136),
.SCD(net125),
.SCE(out46),
.CLK(clk),
.Q(net137)
);

sky130_fd_sc_hd__or4bb_1 c215(
.A(net118),
.B(net67),
.C_N(net129),
.D_N(net134),
.X(net138)
);

sky130_fd_sc_hd__or3_1 c216(
.A(net130),
.B(in22),
.C(net129),
.X(net139)
);

sky130_fd_sc_hd__mux4_1 c217(
.A0(net132),
.A1(net109),
.A2(net139),
.A3(net138),
.S0(net136),
.S1(net128),
.X(net140)
);

sky130_fd_sc_hd__or4bb_2 c218(
.A(net140),
.B(net136),
.C_N(net138),
.D_N(out43),
.X(net141)
);

sky130_fd_sc_hd__nor3_2 c219(
.A(net139),
.B(out11),
.C(net134),
.Y(net142)
);

sky130_fd_sc_hd__and2b_4 c220(
.A_N(net127),
.B(net39),
.X(net143)
);

sky130_fd_sc_hd__nand2b_1 c221(
.A_N(net22),
.B(in59),
.Y(net144)
);

sky130_fd_sc_hd__nor2_2 c222(
.A(in33),
.B(net124),
.Y(net145)
);

sky130_fd_sc_hd__a2111oi_4 c223(
.A1(net72),
.A2(net128),
.B1(net20),
.C1(net135),
.D1(out22),
.Y(net146)
);

sky130_fd_sc_hd__nor2b_4 c224(
.A(net137),
.B_N(net29),
.Y(net147)
);

sky130_fd_sc_hd__and2b_1 c225(
.A_N(in43),
.B(net147),
.X(net148)
);

sky130_fd_sc_hd__and2_1 c226(
.A(net42),
.B(net142),
.X(net149)
);

sky130_fd_sc_hd__and3b_1 c227(
.A_N(net149),
.B(net148),
.C(net114),
.X(net150)
);

sky130_fd_sc_hd__nor2b_4 c228(
.A(net147),
.B_N(net146),
.Y(net151)
);

sky130_fd_sc_hd__nand2b_1 c229(
.A_N(net67),
.B(net85),
.Y(net152)
);

sky130_fd_sc_hd__clkinv_8 c230(
.A(net611),
.Y(net153)
);

sky130_fd_sc_hd__nand2_2 c231(
.A(net149),
.B(net146),
.Y(out8)
);

sky130_fd_sc_hd__nor2b_1 c232(
.A(net151),
.B_N(net152),
.Y(net154)
);

sky130_fd_sc_hd__and3_1 c233(
.A(net25),
.B(out43),
.C(net151),
.X(net155)
);

sky130_fd_sc_hd__dlygate4sd1_1 c234(
.A(net610),
.X(net156)
);

sky130_fd_sc_hd__sdfrbp_2 c235(
.D(net156),
.RESET_B(net121),
.SCD(out8),
.SCE(net128),
.CLK(clk),
.Q(net157)
);

sky130_fd_sc_hd__or2_4 c236(
.A(net154),
.B(net146),
.X(net158)
);

sky130_fd_sc_hd__nor3b_2 c237(
.A(net134),
.B(net151),
.C_N(net156),
.Y(net159)
);

sky130_fd_sc_hd__or4bb_1 c238(
.A(net157),
.B(net20),
.C_N(net156),
.D_N(net152),
.X(net160)
);

sky130_fd_sc_hd__sdfbbn_1 c239(
.D(net124),
.RESET_B(net156),
.SCD(net158),
.SCE(net152),
.SET_B(net160),
.CLK_N(clk),
.Q(net162),
.Q_N(net161)
);

sky130_fd_sc_hd__mux4_1 c240(
.A0(net145),
.A1(net160),
.A2(net143),
.A3(net147),
.S0(out8),
.S1(net152),
.X(net163)
);

sky130_fd_sc_hd__and2_0 c241(
.A(net162),
.B(net657),
.X(net164)
);

sky130_fd_sc_hd__inv_16 c242(
.A(net617),
.Y(net165)
);

sky130_fd_sc_hd__and2b_4 c243(
.A_N(net159),
.B(out0),
.X(net166)
);

sky130_fd_sc_hd__and3_1 c244(
.A(net55),
.B(net20),
.C(net159),
.X(net167)
);

sky130_fd_sc_hd__nand2_1 c245(
.A(net20),
.B(net57),
.Y(out47)
);

sky130_fd_sc_hd__and3_2 c246(
.A(net31),
.B(net144),
.C(out28),
.X(net168)
);

sky130_fd_sc_hd__nand2b_2 c247(
.A_N(net164),
.B(net56),
.Y(out59)
);

sky130_fd_sc_hd__and2b_2 c248(
.A_N(net56),
.B(net49),
.X(net169)
);

sky130_fd_sc_hd__and2_2 c249(
.A(net169),
.B(net114),
.X(out38)
);

sky130_fd_sc_hd__nand3b_4 c250(
.A_N(net142),
.B(out56),
.C(net57),
.Y(net170)
);

sky130_fd_sc_hd__sdfrtn_1 c251(
.D(net166),
.RESET_B(net55),
.SCD(out23),
.SCE(net160),
.CLK_N(clk),
.Q(net171)
);

sky130_fd_sc_hd__and2_2 c252(
.A(in21),
.B(out54),
.X(net172)
);

sky130_fd_sc_hd__nand3_1 c253(
.A(net160),
.B(net172),
.C(net168),
.Y(net173)
);

sky130_fd_sc_hd__or4bb_1 c254(
.A(net170),
.B(out53),
.C_N(net49),
.D_N(out59),
.X(net174)
);

sky130_fd_sc_hd__buf_1 c255(
.A(net617),
.X(net175)
);

sky130_fd_sc_hd__buf_2 c256(
.A(net694),
.X(net176)
);

sky130_fd_sc_hd__sdfbbn_2 c257(
.D(net173),
.RESET_B(net171),
.SCD(out31),
.SCE(out28),
.SET_B(out1),
.CLK_N(clk),
.Q(net178),
.Q_N(net177)
);

sky130_fd_sc_hd__inv_16 c258(
.A(net694),
.Y(out42)
);

sky130_fd_sc_hd__buf_2 c259(
.A(net688),
.X(out50)
);

sky130_fd_sc_hd__nand3b_4 c260(
.A_N(in33),
.B(net178),
.C(net57),
.Y(out18)
);

sky130_fd_sc_hd__a2111o_1 c261(
.A1(net168),
.A2(net172),
.B1(net175),
.C1(net178),
.D1(out53),
.X(net179)
);

sky130_fd_sc_hd__nand3_1 c262(
.A(net144),
.B(net175),
.C(in32),
.Y(out44)
);

sky130_fd_sc_hd__mux4_1 c263(
.A0(net176),
.A1(net172),
.A2(out1),
.A3(net164),
.S0(net168),
.S1(out44),
.X(net180)
);

sky130_fd_sc_hd__and2b_2 c264(
.A_N(net70),
.B(net59),
.X(net181)
);

sky130_fd_sc_hd__nor2_4 c265(
.A(in19),
.B(net70),
.Y(net182)
);

sky130_fd_sc_hd__and2b_4 c266(
.A_N(net181),
.B(in4),
.X(net183)
);

sky130_fd_sc_hd__nor2_2 c267(
.A(in8),
.B(net79),
.Y(net184)
);

sky130_fd_sc_hd__nor2_1 c268(
.A(net74),
.B(net183),
.Y(net185)
);

sky130_fd_sc_hd__and2b_1 c269(
.A_N(in9),
.B(in5),
.X(net186)
);

sky130_fd_sc_hd__or2b_4 c270(
.A(net184),
.B_N(net181),
.X(net187)
);

sky130_fd_sc_hd__nor2_2 c271(
.A(net183),
.B(in15),
.Y(net188)
);

sky130_fd_sc_hd__or2_4 c272(
.A(net64),
.B(in0),
.X(net189)
);

sky130_fd_sc_hd__nand2b_1 c273(
.A_N(in18),
.B(net188),
.Y(net190)
);

sky130_fd_sc_hd__nor2b_2 c274(
.A(in0),
.B_N(net185),
.Y(net191)
);

sky130_fd_sc_hd__nand2_4 c275(
.A(in11),
.B(net184),
.Y(net192)
);

sky130_fd_sc_hd__nand2b_4 c276(
.A_N(net63),
.B(net192),
.Y(net193)
);

sky130_fd_sc_hd__nor2b_4 c277(
.A(net186),
.B_N(net181),
.Y(net194)
);

sky130_fd_sc_hd__nand2b_2 c278(
.A_N(net191),
.B(net184),
.Y(net195)
);

sky130_fd_sc_hd__and3b_2 c279(
.A_N(net191),
.B(net60),
.C(net192),
.X(net196)
);

sky130_fd_sc_hd__nand2_1 c280(
.A(net194),
.B(net182),
.Y(net197)
);

sky130_fd_sc_hd__and2_4 c281(
.A(net195),
.B(net192),
.X(net198)
);

sky130_fd_sc_hd__and3_1 c282(
.A(net189),
.B(net198),
.C(net197),
.X(net199)
);

sky130_fd_sc_hd__nor3_1 c283(
.A(net197),
.B(net199),
.C(net195),
.Y(net200)
);

sky130_fd_sc_hd__or3b_2 c284(
.A(net190),
.B(net200),
.C_N(net197),
.X(net201)
);

sky130_fd_sc_hd__mux4_1 c285(
.A0(net201),
.A1(net195),
.A2(net200),
.A3(net199),
.S0(net193),
.S1(net198),
.X(net202)
);

sky130_fd_sc_hd__nand2_1 c286(
.A(in6),
.B(net88),
.Y(net203)
);

sky130_fd_sc_hd__or2b_1 c287(
.A(in4),
.B_N(net64),
.X(net204)
);

sky130_fd_sc_hd__or2b_2 c288(
.A(net96),
.B_N(net93),
.X(net205)
);

sky130_fd_sc_hd__nand2_2 c289(
.A(net92),
.B(net88),
.Y(net206)
);

sky130_fd_sc_hd__and2_1 c290(
.A(net200),
.B(in10),
.X(net207)
);

sky130_fd_sc_hd__nand2b_4 c291(
.A_N(net206),
.B(net199),
.Y(net208)
);

sky130_fd_sc_hd__nand2_1 c292(
.A(in4),
.B(in29),
.Y(net209)
);

sky130_fd_sc_hd__nor2b_2 c293(
.A(net83),
.B_N(net93),
.Y(net210)
);

sky130_fd_sc_hd__or2_1 c294(
.A(net208),
.B(net209),
.X(net211)
);

sky130_fd_sc_hd__and2_2 c295(
.A(in12),
.B(net96),
.X(net212)
);

sky130_fd_sc_hd__or2b_1 c296(
.A(net203),
.B_N(net210),
.X(net213)
);

sky130_fd_sc_hd__or2_2 c297(
.A(net199),
.B(net213),
.X(net214)
);

sky130_fd_sc_hd__nand2b_2 c298(
.A_N(net210),
.B(net100),
.Y(net215)
);

sky130_fd_sc_hd__or2b_4 c299(
.A(net215),
.B_N(net208),
.X(net216)
);

sky130_fd_sc_hd__nand2b_4 c300(
.A_N(net100),
.B(net206),
.Y(net217)
);

sky130_fd_sc_hd__clkbuf_1 c301(
.A(net684),
.X(net218)
);

sky130_fd_sc_hd__and2b_2 c302(
.A_N(net214),
.B(net205),
.X(net219)
);

sky130_fd_sc_hd__buf_1 c303(
.A(net683),
.X(net220)
);

sky130_fd_sc_hd__nor2_1 c304(
.A(net220),
.B(net217),
.Y(net221)
);

sky130_fd_sc_hd__sdfbbp_1 c305(
.D(net80),
.RESET_B(net221),
.SCD(net88),
.SCE(net220),
.SET_B(net211),
.CLK(clk),
.Q(net223),
.Q_N(net222)
);

sky130_fd_sc_hd__nand2_2 c306(
.A(net188),
.B(net220),
.Y(net224)
);

sky130_fd_sc_hd__sdfbbn_1 c307(
.D(net224),
.RESET_B(in41),
.SCD(net219),
.SCE(net220),
.SET_B(net195),
.CLK_N(clk),
.Q(net225)
);

sky130_fd_sc_hd__nor2b_4 c308(
.A(net122),
.B_N(net205),
.Y(net226)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c309(
.A(net630),
.X(net227)
);

sky130_fd_sc_hd__and2b_2 c310(
.A_N(net97),
.B(net116),
.X(net228)
);

sky130_fd_sc_hd__nand2b_1 c311(
.A_N(net206),
.B(in58),
.Y(net229)
);

sky130_fd_sc_hd__inv_12 c312(
.A(net631),
.Y(net230)
);

sky130_fd_sc_hd__nor2_1 c313(
.A(net229),
.B(net230),
.Y(net231)
);

sky130_fd_sc_hd__nor3b_2 c314(
.A(in17),
.B(in21),
.C_N(net230),
.Y(net232)
);

sky130_fd_sc_hd__or2b_1 c315(
.A(net197),
.B_N(net229),
.X(net233)
);

sky130_fd_sc_hd__or3b_2 c316(
.A(net233),
.B(net231),
.C_N(net193),
.X(net234)
);

sky130_fd_sc_hd__and2_0 c317(
.A(net231),
.B(out52),
.X(net235)
);

sky130_fd_sc_hd__nand2b_4 c318(
.A_N(net230),
.B(net189),
.Y(net236)
);

sky130_fd_sc_hd__or3b_4 c319(
.A(net236),
.B(net122),
.C_N(net85),
.X(net237)
);

sky130_fd_sc_hd__and2b_4 c320(
.A_N(net107),
.B(net229),
.X(net238)
);

sky130_fd_sc_hd__nor2_2 c321(
.A(net238),
.B(in34),
.Y(net239)
);

sky130_fd_sc_hd__and2_4 c322(
.A(net71),
.B(net183),
.X(net240)
);

sky130_fd_sc_hd__and3b_4 c323(
.A_N(net235),
.B(net230),
.C(net71),
.X(net241)
);

sky130_fd_sc_hd__nand2_4 c324(
.A(net209),
.B(net231),
.Y(net242)
);

sky130_fd_sc_hd__dlygate4sd1_1 c325(
.A(net693),
.X(net243)
);

sky130_fd_sc_hd__mux4_2 c326(
.A0(net239),
.A1(net105),
.A2(net243),
.A3(net228),
.S0(in0),
.S1(net230),
.X(net244)
);

sky130_fd_sc_hd__buf_8 c327(
.A(net692),
.X(out2)
);

sky130_fd_sc_hd__sdfrtp_1 c328(
.D(net240),
.RESET_B(net244),
.SCD(net237),
.SCE(net114),
.CLK(clk),
.Q(net245)
);

sky130_fd_sc_hd__mux4_4 c329(
.A0(net226),
.A1(net229),
.A2(net245),
.A3(net244),
.S0(net241),
.S1(net243),
.X(net246)
);

sky130_fd_sc_hd__a2111o_4 c330(
.A1(net141),
.A2(net59),
.B1(in29),
.C1(net135),
.D1(net245),
.X(net247)
);

sky130_fd_sc_hd__clkbuf_1 c331(
.A(net607),
.X(net248)
);

sky130_fd_sc_hd__and2_2 c332(
.A(net242),
.B(in7),
.X(net249)
);

sky130_fd_sc_hd__nand2_1 c333(
.A(net21),
.B(net244),
.Y(out21)
);

sky130_fd_sc_hd__or2_2 c334(
.A(net138),
.B(net128),
.X(out35)
);

sky130_fd_sc_hd__nand2b_2 c335(
.A_N(net89),
.B(net138),
.Y(net250)
);

sky130_fd_sc_hd__or2b_2 c336(
.A(net131),
.B_N(net89),
.X(net251)
);

sky130_fd_sc_hd__or2_1 c337(
.A(net23),
.B(net121),
.X(net252)
);

sky130_fd_sc_hd__and2b_4 c338(
.A_N(net244),
.B(net252),
.X(out3)
);

sky130_fd_sc_hd__or3_1 c339(
.A(net251),
.B(in49),
.C(net59),
.X(net253)
);

sky130_fd_sc_hd__nor2_2 c340(
.A(net204),
.B(net252),
.Y(net254)
);

sky130_fd_sc_hd__and2b_1 c341(
.A_N(net228),
.B(out43),
.X(net255)
);

sky130_fd_sc_hd__or2b_2 c342(
.A(net252),
.B_N(net184),
.X(net256)
);

sky130_fd_sc_hd__buf_2 c343(
.A(net606),
.X(net257)
);

sky130_fd_sc_hd__nand2_2 c344(
.A(net253),
.B(net659),
.Y(net258)
);

sky130_fd_sc_hd__or2b_4 c345(
.A(net205),
.B_N(net245),
.X(net259)
);

sky130_fd_sc_hd__nor2_1 c346(
.A(net259),
.B(net252),
.Y(net260)
);

sky130_fd_sc_hd__dlygate4sd3_1 c347(
.A(net651),
.X(net261)
);

sky130_fd_sc_hd__clkinv_2 c348(
.A(net651),
.Y(net262)
);

sky130_fd_sc_hd__sdfrtp_2 c349(
.D(net255),
.RESET_B(out11),
.SCD(net119),
.SCE(net254),
.CLK(clk),
.Q(net263)
);

sky130_fd_sc_hd__sdfbbn_2 c350(
.D(net258),
.RESET_B(net204),
.SCD(net4),
.SCE(net254),
.SET_B(net256),
.CLK_N(clk),
.Q(net265),
.Q_N(net264)
);

sky130_fd_sc_hd__and2b_1 c351(
.A_N(net257),
.B(net23),
.X(out25)
);

sky130_fd_sc_hd__nor3_2 c352(
.A(net187),
.B(net85),
.C(in53),
.Y(out45)
);

sky130_fd_sc_hd__inv_8 c353(
.A(net608),
.Y(out6)
);

sky130_fd_sc_hd__sdfrtp_4 c354(
.D(net253),
.RESET_B(net153),
.SCD(net135),
.SCE(net254),
.CLK(clk),
.Q(net266)
);

sky130_fd_sc_hd__buf_2 c355(
.A(net691),
.X(out36)
);

sky130_fd_sc_hd__nor2b_1 c356(
.A(net15),
.B_N(net146),
.Y(net267)
);

sky130_fd_sc_hd__buf_4 c357(
.A(net690),
.X(net268)
);

sky130_fd_sc_hd__o2111ai_2 c358(
.A1(net232),
.A2(in7),
.B1(out22),
.C1(net152),
.D1(net268),
.Y(net269)
);

sky130_fd_sc_hd__dfbbn_1 c359(
.D(net158),
.RESET_B(out56),
.SET_B(net657),
.CLK_N(clk),
.Q(net270)
);

sky130_fd_sc_hd__and2_1 c360(
.A(net234),
.B(net34),
.X(out57)
);

sky130_fd_sc_hd__and2_4 c361(
.A(net155),
.B(net39),
.X(net271)
);

sky130_fd_sc_hd__nor3_4 c362(
.A(net161),
.B(net267),
.C(in53),
.Y(net272)
);

sky130_fd_sc_hd__dfbbn_2 c363(
.D(in59),
.RESET_B(out45),
.SET_B(out57),
.CLK_N(clk),
.Q(out60),
.Q_N(net273)
);

sky130_fd_sc_hd__or3_2 c364(
.A(net152),
.B(net2),
.C(net273),
.X(out16)
);

sky130_fd_sc_hd__dfbbp_1 c365(
.D(net271),
.RESET_B(net155),
.SET_B(net267),
.CLK(clk),
.Q(net275),
.Q_N(net274)
);

sky130_fd_sc_hd__and3b_4 c366(
.A_N(net269),
.B(out45),
.C(net250),
.X(net276)
);

sky130_fd_sc_hd__nand3b_1 c367(
.A_N(net250),
.B(out16),
.C(net34),
.Y(net277)
);

sky130_fd_sc_hd__or3b_2 c368(
.A(net135),
.B(net268),
.C_N(net272),
.X(out49)
);

sky130_fd_sc_hd__or3b_2 c369(
.A(net99),
.B(net274),
.C_N(net276),
.X(net278)
);

sky130_fd_sc_hd__and2_0 c370(
.A(net245),
.B(net275),
.X(net279)
);

sky130_fd_sc_hd__inv_16 c371(
.A(net695),
.Y(out58)
);

sky130_fd_sc_hd__dlygate4sd3_1 c372(
.A(net609),
.X(out55)
);

sky130_fd_sc_hd__mux4_4 c373(
.A0(net270),
.A1(net268),
.A2(net253),
.A3(net187),
.S0(net146),
.S1(net276),
.X(net280)
);

sky130_fd_sc_hd__mux4_1 c392(
.A0(net179),
.A1(in43),
.A2(out25),
.A3(out43),
.S0(out2),
.S1(out53),
.X(net281)
);

sky130_fd_sc_hd__sdfbbp_1 c393(
.D(net58),
.RESET_B(out43),
.SCD(out8),
.SCE(out31),
.SET_B(out24),
.CLK(clk),
.Q(out30)
);

sky130_fd_sc_hd__mux4_2 c394(
.A0(net165),
.A1(net279),
.A2(net59),
.A3(out44),
.S0(out54),
.S1(out24),
.X(out51)
);

sky130_fd_sc_hd__mux4_2 c395(
.A0(net49),
.A1(net121),
.A2(out2),
.A3(out8),
.S0(net658),
.S1(out24),
.X(net282)
);

sky130_fd_sc_hd__or4bb_4 c396(
.A(in1),
.B(net188),
.C_N(in0),
.D_N(net198),
.X(net283)
);

sky130_fd_sc_hd__nand2b_4 c397(
.A_N(in14),
.B(net185),
.Y(net284)
);

sky130_fd_sc_hd__or2b_2 c398(
.A(net193),
.B_N(net77),
.X(net285)
);

sky130_fd_sc_hd__or2_2 c399(
.A(net285),
.B(net198),
.X(net286)
);

sky130_fd_sc_hd__or2_2 c400(
.A(net286),
.B(net193),
.X(net287)
);

sky130_fd_sc_hd__and2_0 c401(
.A(net196),
.B(net64),
.X(net288)
);

sky130_fd_sc_hd__nand2b_4 c402(
.A_N(net188),
.B(net284),
.Y(net289)
);

sky130_fd_sc_hd__nor2_4 c403(
.A(net182),
.B(net185),
.Y(net290)
);

sky130_fd_sc_hd__and2_2 c404(
.A(net288),
.B(net289),
.X(net291)
);

sky130_fd_sc_hd__and2_2 c405(
.A(net290),
.B(net79),
.X(net292)
);

sky130_fd_sc_hd__or2_2 c406(
.A(net185),
.B(net286),
.X(net293)
);

sky130_fd_sc_hd__nor2b_4 c407(
.A(net288),
.B_N(net291),
.Y(net294)
);

sky130_fd_sc_hd__clkinv_4 c408(
.A(net644),
.Y(net295)
);

sky130_fd_sc_hd__nand2b_2 c409(
.A_N(net192),
.B(net288),
.Y(net296)
);

sky130_fd_sc_hd__nand2_2 c410(
.A(net190),
.B(net290),
.Y(net297)
);

sky130_fd_sc_hd__sdfbbn_1 c411(
.D(net297),
.RESET_B(net295),
.SCD(net285),
.SCE(net287),
.SET_B(net291),
.CLK_N(clk),
.Q(net299),
.Q_N(net298)
);

sky130_fd_sc_hd__nand2_1 c412(
.A(net194),
.B(net192),
.Y(net300)
);

sky130_fd_sc_hd__or2b_1 c413(
.A(net300),
.B_N(net77),
.X(net301)
);

sky130_fd_sc_hd__and2_2 c414(
.A(net291),
.B(net290),
.X(net302)
);

sky130_fd_sc_hd__and2b_2 c415(
.A_N(in14),
.B(net300),
.X(net303)
);

sky130_fd_sc_hd__nand2b_2 c416(
.A_N(net303),
.B(net297),
.Y(net304)
);

sky130_fd_sc_hd__mux4_4 c417(
.A0(net289),
.A1(net293),
.A2(net304),
.A3(net292),
.S0(net291),
.S1(net294),
.X(net305)
);

sky130_fd_sc_hd__and2b_2 c418(
.A_N(net220),
.B(in23),
.X(net306)
);

sky130_fd_sc_hd__nand3_4 c419(
.A(net300),
.B(net77),
.C(net284),
.Y(net307)
);

sky130_fd_sc_hd__or2b_4 c420(
.A(net215),
.B_N(net285),
.X(net308)
);

sky130_fd_sc_hd__sdfxbp_1 c421(
.D(net186),
.SCD(net308),
.SCE(net220),
.CLK(clk),
.Q(net309)
);

sky130_fd_sc_hd__nor3_4 c422(
.A(net297),
.B(net307),
.C(net291),
.Y(net310)
);

sky130_fd_sc_hd__and3_1 c423(
.A(net225),
.B(in17),
.C(net184),
.X(net311)
);

sky130_fd_sc_hd__inv_2 c424(
.A(net624),
.Y(net312)
);

sky130_fd_sc_hd__and3_1 c425(
.A(net224),
.B(net283),
.C(net284),
.X(net313)
);

sky130_fd_sc_hd__nor2_2 c426(
.A(net313),
.B(in23),
.Y(net314)
);

sky130_fd_sc_hd__nand3_2 c427(
.A(net312),
.B(net212),
.C(net298),
.Y(net315)
);

sky130_fd_sc_hd__sdfxbp_2 c428(
.D(in35),
.SCD(net308),
.SCE(net292),
.CLK(clk),
.Q(net317),
.Q_N(net316)
);

sky130_fd_sc_hd__buf_4 c429(
.A(net623),
.X(net318)
);

sky130_fd_sc_hd__or3_1 c430(
.A(net283),
.B(net313),
.C(net312),
.X(net319)
);

sky130_fd_sc_hd__clkbuf_4 c431(
.A(net644),
.X(net320)
);

sky130_fd_sc_hd__or3b_2 c432(
.A(net309),
.B(net318),
.C_N(net312),
.X(net321)
);

sky130_fd_sc_hd__sdfxtp_1 c433(
.D(net311),
.SCD(net314),
.SCE(net306),
.CLK(clk),
.Q(net322)
);

sky130_fd_sc_hd__nor2b_1 c434(
.A(net321),
.B_N(net320),
.Y(net323)
);

sky130_fd_sc_hd__and3b_2 c435(
.A_N(net212),
.B(net320),
.C(net322),
.X(net324)
);

sky130_fd_sc_hd__mux4_2 c436(
.A0(net323),
.A1(net312),
.A2(net324),
.A3(net284),
.S0(net216),
.S1(net314),
.X(net325)
);

sky130_fd_sc_hd__mux4_1 c437(
.A0(net322),
.A1(net317),
.A2(net315),
.A3(net318),
.S0(net213),
.S1(net220),
.X(net326)
);

sky130_fd_sc_hd__mux4_2 c438(
.A0(net326),
.A1(net324),
.A2(net313),
.A3(net287),
.S0(net292),
.S1(net661),
.X(net327)
);

sky130_fd_sc_hd__sdfbbn_2 c439(
.D(net302),
.RESET_B(net326),
.SCD(net186),
.SCE(net215),
.SET_B(net662),
.CLK_N(clk),
.Q(net328)
);

sky130_fd_sc_hd__or3b_2 c440(
.A(net203),
.B(net227),
.C_N(net663),
.X(net329)
);

sky130_fd_sc_hd__nor3_2 c441(
.A(net189),
.B(net222),
.C(net329),
.Y(out7)
);

sky130_fd_sc_hd__nor3_1 c442(
.A(net208),
.B(net101),
.C(net329),
.Y(net330)
);

sky130_fd_sc_hd__nand3_2 c443(
.A(net101),
.B(net243),
.C(out7),
.Y(net331)
);

sky130_fd_sc_hd__a2111oi_0 c444(
.A1(net304),
.A2(net101),
.B1(net116),
.C1(net243),
.D1(net315),
.Y(net332)
);

sky130_fd_sc_hd__or3_2 c445(
.A(net0),
.B(net227),
.C(out7),
.X(out5)
);

sky130_fd_sc_hd__clkinv_16 c446(
.A(net628),
.Y(net333)
);

sky130_fd_sc_hd__or3b_1 c447(
.A(net102),
.B(net243),
.C_N(net116),
.X(net334)
);

sky130_fd_sc_hd__nand2b_4 c448(
.A_N(net223),
.B(in59),
.Y(net335)
);

sky130_fd_sc_hd__and2b_2 c449(
.A_N(net315),
.B(net296),
.X(net336)
);

sky130_fd_sc_hd__nand2b_2 c450(
.A_N(net227),
.B(net241),
.Y(net337)
);

sky130_fd_sc_hd__or2_4 c451(
.A(net335),
.B(in58),
.X(net338)
);

sky130_fd_sc_hd__nor3b_4 c452(
.A(net285),
.B(out5),
.C_N(out7),
.Y(net339)
);

sky130_fd_sc_hd__inv_6 c453(
.A(net627),
.Y(net340)
);

sky130_fd_sc_hd__sdfsbp_1 c454(
.D(net329),
.SCD(out22),
.SCE(net331),
.SET_B(in58),
.CLK(clk),
.Q(net342),
.Q_N(net341)
);

sky130_fd_sc_hd__or4bb_4 c455(
.A(net328),
.B(net329),
.C_N(net335),
.D_N(net340),
.X(net343)
);

sky130_fd_sc_hd__mux4_1 c456(
.A0(net331),
.A1(net338),
.A2(net340),
.A3(net339),
.S0(net102),
.S1(net336),
.X(net344)
);

sky130_fd_sc_hd__sdfxtp_2 c457(
.D(net319),
.SCD(net227),
.SCE(net340),
.CLK(clk),
.Q(net345)
);

sky130_fd_sc_hd__nand3_1 c458(
.A(net339),
.B(net296),
.C(net333),
.Y(out14)
);

sky130_fd_sc_hd__sdfxtp_4 c459(
.D(net333),
.SCD(net336),
.SCE(net341),
.CLK(clk),
.Q(net346)
);

sky130_fd_sc_hd__mux4_2 c460(
.A0(net346),
.A1(net334),
.A2(net336),
.A3(net241),
.S0(net285),
.S1(net340),
.X(net347)
);

sky130_fd_sc_hd__or4bb_4 c461(
.A(net342),
.B(net345),
.C_N(net346),
.D_N(net666),
.X(net348)
);

sky130_fd_sc_hd__dfbbn_1 c462(
.D(net187),
.RESET_B(net254),
.SET_B(net337),
.CLK_N(clk),
.Q(net350),
.Q_N(net349)
);

sky130_fd_sc_hd__dfbbn_2 c463(
.D(net8),
.RESET_B(net287),
.SET_B(net320),
.CLK_N(clk),
.Q(net351)
);

sky130_fd_sc_hd__or2_1 c464(
.A(net243),
.B(net292),
.X(net352)
);

sky130_fd_sc_hd__nor2b_1 c465(
.A(net307),
.B_N(net340),
.Y(net353)
);

sky130_fd_sc_hd__nor2_4 c466(
.A(net337),
.B(net349),
.Y(net354)
);

sky130_fd_sc_hd__nand2b_4 c467(
.A_N(net340),
.B(net307),
.Y(net355)
);

sky130_fd_sc_hd__nand2b_1 c468(
.A_N(net320),
.B(net352),
.Y(net356)
);

sky130_fd_sc_hd__inv_4 c469(
.A(net613),
.Y(net357)
);

sky130_fd_sc_hd__sdfbbp_1 c470(
.D(net350),
.RESET_B(net262),
.SCD(net324),
.SCE(net308),
.SET_B(out2),
.CLK(clk),
.Q(net358)
);

sky130_fd_sc_hd__or2_4 c471(
.A(net296),
.B(net261),
.X(net359)
);

sky130_fd_sc_hd__buf_6 c472(
.A(net613),
.X(net360)
);

sky130_fd_sc_hd__nor2b_1 c473(
.A(net343),
.B_N(net263),
.Y(net361)
);

sky130_fd_sc_hd__mux4_2 c474(
.A0(net356),
.A1(net18),
.A2(net316),
.A3(out2),
.S0(net357),
.S1(net119),
.X(net362)
);

sky130_fd_sc_hd__nand2b_2 c475(
.A_N(net261),
.B(net352),
.Y(net363)
);

sky130_fd_sc_hd__sdfsbp_2 c476(
.D(net360),
.SCD(net243),
.SCE(net354),
.SET_B(net352),
.CLK(clk),
.Q(out29),
.Q_N(net364)
);

sky130_fd_sc_hd__sdfstp_1 c477(
.D(net287),
.SCD(net361),
.SCE(net364),
.SET_B(net256),
.CLK(clk),
.Q(net365)
);

sky130_fd_sc_hd__sdfbbn_1 c478(
.D(net248),
.RESET_B(net265),
.SCD(net343),
.SCE(net354),
.SET_B(net316),
.CLK_N(clk),
.Q(net367),
.Q_N(net366)
);

sky130_fd_sc_hd__o2111a_2 c479(
.A1(net367),
.A2(net364),
.B1(net340),
.C1(net248),
.D1(in53),
.X(out33)
);

sky130_fd_sc_hd__or3b_1 c480(
.A(net355),
.B(net357),
.C_N(in21),
.X(net368)
);

sky130_fd_sc_hd__dfbbp_1 c481(
.D(net354),
.RESET_B(out29),
.SET_B(out33),
.CLK(clk),
.Q(net369)
);

sky130_fd_sc_hd__nand3_4 c482(
.A(net184),
.B(net369),
.C(net193),
.Y(net370)
);

sky130_fd_sc_hd__sdfbbn_2 c483(
.D(net363),
.RESET_B(net366),
.SCD(net368),
.SCE(out33),
.SET_B(net365),
.CLK_N(clk),
.Q(net371)
);

sky130_fd_sc_hd__and2_4 c484(
.A(net121),
.B(net668),
.X(net372)
);

sky130_fd_sc_hd__nor3_1 c485(
.A(net2),
.B(net324),
.C(net266),
.Y(net373)
);

sky130_fd_sc_hd__nand3_2 c486(
.A(net312),
.B(net4),
.C(out7),
.Y(net374)
);

sky130_fd_sc_hd__or2b_4 c487(
.A(net267),
.B_N(net273),
.X(net375)
);

sky130_fd_sc_hd__inv_12 c488(
.A(net688),
.Y(net376)
);

sky130_fd_sc_hd__buf_8 c489(
.X(net377)
);

sky130_fd_sc_hd__sdfstp_2 c490(
.D(net371),
.SCD(out8),
.SCE(out33),
.SET_B(out7),
.CLK(clk),
.Q(out37)
);

sky130_fd_sc_hd__or3_1 c491(
.A(net374),
.B(net241),
.C(net665),
.X(net378)
);

sky130_fd_sc_hd__dlygate4sd3_1 c492(
.A(net689),
.X(out10)
);

sky130_fd_sc_hd__inv_4 c493(
.A(net604),
.Y(net379)
);

sky130_fd_sc_hd__or3_1 c494(
.A(net148),
.B(net267),
.C(net664),
.X(net380)
);

sky130_fd_sc_hd__nand2_4 c495(
.A(net324),
.B(out2),
.Y(out32)
);

sky130_fd_sc_hd__nor3_4 c496(
.A(net153),
.B(out36),
.C(net317),
.Y(net381)
);

sky130_fd_sc_hd__nor3b_2 c497(
.A(net380),
.B(out36),
.C_N(net39),
.Y(net382)
);

sky130_fd_sc_hd__inv_1 c498(
.A(net689),
.Y(net383)
);

sky130_fd_sc_hd__nor3b_1 c499(
.A(net266),
.B(net381),
.C_N(net39),
.Y(net384)
);

sky130_fd_sc_hd__sdfbbp_1 c500(
.D(net59),
.RESET_B(net383),
.SCD(net378),
.SCE(out36),
.SET_B(out3),
.CLK(clk),
.Q(net386),
.Q_N(net385)
);

sky130_fd_sc_hd__nand3_2 c501(
.A(net39),
.B(net377),
.C(net385),
.Y(net387)
);

sky130_fd_sc_hd__and3b_2 c502(
.A_N(net291),
.B(net379),
.C(out33),
.X(net388)
);

sky130_fd_sc_hd__or4bb_2 c503(
.A(net183),
.B(net386),
.C_N(net324),
.D_N(net280),
.X(net389)
);

sky130_fd_sc_hd__sdfstp_4 c504(
.D(net388),
.SCD(net389),
.SCE(net386),
.SET_B(net387),
.CLK(clk),
.Q(out26)
);

sky130_fd_sc_hd__or4bb_2 c505(
.A(net146),
.B(net384),
.C_N(net385),
.D_N(net4),
.X(net390)
);

sky130_fd_sc_hd__and2_2 c528(
.A(net79),
.B(net292),
.X(net391)
);

sky130_fd_sc_hd__nor2b_1 c529(
.A(net295),
.B_N(in21),
.Y(net392)
);

sky130_fd_sc_hd__nor2b_4 c530(
.A(net60),
.B_N(net295),
.Y(net393)
);

sky130_fd_sc_hd__nor2_2 c531(
.A(net283),
.B(net392),
.Y(net394)
);

sky130_fd_sc_hd__and2_4 c532(
.A(net286),
.B(net196),
.X(net395)
);

sky130_fd_sc_hd__and2b_1 c533(
.A_N(net392),
.B(net391),
.X(net396)
);

sky130_fd_sc_hd__clkbuf_1 c534(
.X(net397)
);

sky130_fd_sc_hd__clkinv_2 c535(
.A(net632),
.Y(net398)
);

sky130_fd_sc_hd__inv_1 c536(
.A(net653),
.Y(net399)
);

sky130_fd_sc_hd__clkinv_2 c537(
.A(net653),
.Y(net400)
);

sky130_fd_sc_hd__nor2_4 c538(
.A(net394),
.B(net392),
.Y(net401)
);

sky130_fd_sc_hd__dfrbp_1 c539(
.D(net395),
.RESET_B(net399),
.CLK(clk),
.Q(net402)
);

sky130_fd_sc_hd__or2_1 c540(
.A(net400),
.B(net391),
.X(net403)
);

sky130_fd_sc_hd__nand2_4 c541(
.A(net396),
.B(net397),
.Y(net404)
);

sky130_fd_sc_hd__nor2b_1 c542(
.A(net399),
.B_N(net660),
.Y(net405)
);

sky130_fd_sc_hd__or2b_4 c543(
.A(net398),
.B_N(net405),
.X(net406)
);

sky130_fd_sc_hd__nor2b_4 c544(
.A(net402),
.B_N(net406),
.Y(net407)
);

sky130_fd_sc_hd__nand2b_1 c545(
.A_N(net405),
.B(net195),
.Y(net408)
);

sky130_fd_sc_hd__dfrbp_2 c546(
.D(net401),
.RESET_B(net400),
.CLK(clk),
.Q(net410),
.Q_N(net409)
);

sky130_fd_sc_hd__or2b_4 c547(
.A(net407),
.B_N(net408),
.X(net411)
);

sky130_fd_sc_hd__and2_2 c548(
.A(net408),
.B(net405),
.X(net412)
);

sky130_fd_sc_hd__nand2b_1 c549(
.A_N(net404),
.B(net408),
.Y(net413)
);

sky130_fd_sc_hd__nand2b_2 c550(
.A_N(in17),
.B(net93),
.Y(net414)
);

sky130_fd_sc_hd__or2_1 c551(
.A(in23),
.B(net195),
.X(net415)
);

sky130_fd_sc_hd__inv_2 c552(
.A(net633),
.Y(net416)
);

sky130_fd_sc_hd__and2_2 c553(
.A(net406),
.B(net660),
.X(net417)
);

sky130_fd_sc_hd__and2_1 c554(
.A(net415),
.B(net306),
.X(net418)
);

sky130_fd_sc_hd__or2b_1 c555(
.A(in1),
.B_N(net660),
.X(net419)
);

sky130_fd_sc_hd__or2b_4 c556(
.A(net213),
.B_N(net79),
.X(net420)
);

sky130_fd_sc_hd__nor2_1 c557(
.A(net195),
.B(net410),
.Y(net421)
);

sky130_fd_sc_hd__nand2_2 c558(
.A(net77),
.B(net217),
.Y(net422)
);

sky130_fd_sc_hd__buf_6 c559(
.A(net633),
.X(net423)
);

sky130_fd_sc_hd__and2_0 c560(
.A(net418),
.B(net391),
.X(net424)
);

sky130_fd_sc_hd__and2_2 c561(
.A(net417),
.B(net661),
.X(net425)
);

sky130_fd_sc_hd__nand3b_4 c562(
.A_N(net420),
.B(net410),
.C(net424),
.Y(net426)
);

sky130_fd_sc_hd__dfrtn_1 c563(
.D(net414),
.RESET_B(net319),
.CLK_N(clk),
.Q(net427)
);

sky130_fd_sc_hd__and2b_1 c564(
.A_N(net421),
.B(net411),
.X(net428)
);

sky130_fd_sc_hd__a2111oi_1 c565(
.A1(net419),
.A2(net198),
.B1(net424),
.C1(net423),
.D1(net316),
.Y(net429)
);

sky130_fd_sc_hd__o2111a_4 c566(
.A1(net306),
.A2(net299),
.B1(net318),
.C1(net415),
.D1(net424),
.X(net430)
);

sky130_fd_sc_hd__buf_1 c567(
.A(net642),
.X(net431)
);

sky130_fd_sc_hd__sdfbbn_1 c568(
.D(net423),
.RESET_B(net284),
.SCD(net431),
.SCE(net424),
.SET_B(net314),
.CLK_N(clk),
.Q(net433),
.Q_N(net432)
);

sky130_fd_sc_hd__sedfxbp_1 c569(
.D(net429),
.DE(net430),
.SCD(net432),
.SCE(net424),
.CLK(clk),
.Q(net434)
);

sky130_fd_sc_hd__dfrtp_1 c570(
.D(net426),
.RESET_B(in5),
.CLK(clk),
.Q(net435)
);

sky130_fd_sc_hd__or4bb_4 c571(
.A(net434),
.B(net433),
.C_N(net435),
.D_N(net424),
.X(net436)
);

sky130_fd_sc_hd__and2_1 c572(
.A(net318),
.B(net93),
.X(net437)
);

sky130_fd_sc_hd__clkinv_16 c573(
.A(net612),
.Y(net438)
);

sky130_fd_sc_hd__and2b_4 c574(
.A_N(net437),
.B(net663),
.X(net439)
);

sky130_fd_sc_hd__nand2_1 c575(
.A(net116),
.B(net435),
.Y(net440)
);

sky130_fd_sc_hd__nor3_1 c576(
.A(net416),
.B(net440),
.C(net661),
.Y(net441)
);

sky130_fd_sc_hd__and3_1 c577(
.A(net440),
.B(out7),
.C(net196),
.X(net442)
);

sky130_fd_sc_hd__sdfbbn_2 c578(
.D(net105),
.RESET_B(net437),
.SCD(net336),
.SCE(net114),
.SET_B(net663),
.CLK_N(clk),
.Q(net443)
);

sky130_fd_sc_hd__and3_2 c579(
.A(net442),
.B(net241),
.C(net440),
.X(net444)
);

sky130_fd_sc_hd__nand2b_4 c580(
.A_N(net444),
.B(net318),
.Y(net445)
);

sky130_fd_sc_hd__buf_2 c581(
.A(net612),
.X(net446)
);

sky130_fd_sc_hd__inv_16 c582(
.A(net643),
.Y(net447)
);

sky130_fd_sc_hd__or3b_1 c583(
.A(net411),
.B(net440),
.C_N(net406),
.X(net448)
);

sky130_fd_sc_hd__buf_4 c584(
.A(net646),
.X(net449)
);

sky130_fd_sc_hd__sdfxbp_1 c585(
.D(net445),
.SCD(net443),
.SCE(net449),
.CLK(clk),
.Q(net450)
);

sky130_fd_sc_hd__dlymetal6s2s_1 c586(
.A(net655),
.X(net451)
);

sky130_fd_sc_hd__and2_0 c587(
.A(net439),
.B(net449),
.X(net452)
);

sky130_fd_sc_hd__or3_1 c588(
.A(net447),
.B(net451),
.C(net667),
.X(net453)
);

sky130_fd_sc_hd__sdfbbp_1 c589(
.D(net406),
.RESET_B(net123),
.SCD(net336),
.SCE(in59),
.SET_B(net292),
.CLK(clk),
.Q(net455),
.Q_N(net454)
);

sky130_fd_sc_hd__mux4_1 c590(
.A0(net447),
.A1(net455),
.A2(net440),
.A3(net453),
.S0(net424),
.S1(net451),
.X(net456)
);

sky130_fd_sc_hd__o2111a_4 c591(
.A1(net452),
.A2(net241),
.B1(net453),
.C1(net454),
.D1(net661),
.X(net457)
);

sky130_fd_sc_hd__mux4_1 c592(
.A0(net456),
.A1(in21),
.A2(net455),
.A3(net348),
.S0(net451),
.S1(net457),
.X(net458)
);

sky130_fd_sc_hd__mux4_4 c593(
.A0(net451),
.A1(net454),
.A2(net440),
.A3(net424),
.S0(net446),
.S1(net669),
.X(net459)
);

sky130_fd_sc_hd__or3_4 c594(
.A(net136),
.B(out2),
.C(net393),
.X(out9)
);

sky130_fd_sc_hd__and2_2 c595(
.A(net334),
.B(net424),
.X(net460)
);

sky130_fd_sc_hd__sdfxbp_2 c596(
.D(net441),
.SCD(net299),
.SCE(out21),
.CLK(clk),
.Q(net462),
.Q_N(net461)
);

sky130_fd_sc_hd__buf_6 c597(
.A(net629),
.X(net463)
);

sky130_fd_sc_hd__nand2_1 c598(
.A(net289),
.B(net193),
.Y(net464)
);

sky130_fd_sc_hd__or3b_4 c599(
.A(net464),
.B(net461),
.C_N(net457),
.X(net465)
);

sky130_fd_sc_hd__sdfxtp_1 c600(
.D(net193),
.SCD(net136),
.SCE(net465),
.CLK(clk),
.Q(net466)
);

sky130_fd_sc_hd__and2b_4 c601(
.A_N(net466),
.B(in15),
.X(out19)
);

sky130_fd_sc_hd__clkinv_1 c602(
.A(net629),
.Y(net467)
);

sky130_fd_sc_hd__buf_2 c603(
.A(net656),
.X(net468)
);

sky130_fd_sc_hd__and2b_2 c604(
.A_N(net353),
.B(net351),
.X(net469)
);

sky130_fd_sc_hd__sdfbbn_1 c605(
.D(net462),
.RESET_B(out3),
.SCD(net465),
.SCE(net306),
.SET_B(net467),
.CLK_N(clk),
.Q(net471),
.Q_N(net470)
);

sky130_fd_sc_hd__o2111ai_1 c606(
.A1(net467),
.A2(net317),
.B1(net457),
.C1(net470),
.D1(net193),
.Y(out13)
);

sky130_fd_sc_hd__sdfxtp_2 c607(
.D(net256),
.SCD(net435),
.SCE(net467),
.CLK(clk),
.Q(net472)
);

sky130_fd_sc_hd__sdfxtp_4 c608(
.D(net336),
.SCD(net370),
.SCE(net393),
.CLK(clk),
.Q(net473)
);

sky130_fd_sc_hd__mux4_1 c609(
.A0(net460),
.A1(net471),
.A2(net301),
.A3(net292),
.S0(net463),
.S1(out19),
.X(net474)
);

sky130_fd_sc_hd__nand3_4 c610(
.A(net472),
.B(net468),
.C(out2),
.Y(net475)
);

sky130_fd_sc_hd__and3_1 c611(
.A(net475),
.B(net467),
.C(net471),
.X(net476)
);

sky130_fd_sc_hd__clkinv_8 c612(
.A(net646),
.Y(out20)
);

sky130_fd_sc_hd__or2b_1 c613(
.A(net18),
.B_N(net467),
.X(net477)
);

sky130_fd_sc_hd__dfbbn_1 c614(
.D(net119),
.RESET_B(net348),
.SET_B(out22),
.CLK_N(clk),
.Q(net478)
);

sky130_fd_sc_hd__sdfbbn_2 c615(
.D(net473),
.RESET_B(net465),
.SCD(net471),
.SCE(net352),
.SET_B(net467),
.CLK_N(clk),
.Q(net479)
);

sky130_fd_sc_hd__or4bb_1 c616(
.A(net438),
.B(net278),
.C_N(out11),
.D_N(net298),
.X(net480)
);

sky130_fd_sc_hd__nor3b_2 c617(
.A(in32),
.B(net306),
.C_N(net299),
.Y(net481)
);

sky130_fd_sc_hd__and3b_1 c618(
.A_N(in15),
.B(net365),
.C(net44),
.X(net482)
);

sky130_fd_sc_hd__and3b_4 c619(
.A_N(net128),
.B(out60),
.C(net241),
.X(out15)
);

sky130_fd_sc_hd__clkbuf_16 c620(
.A(net685),
.X(net483)
);

sky130_fd_sc_hd__and3b_1 c621(
.A_N(in49),
.B(net123),
.C(out22),
.X(net484)
);

sky130_fd_sc_hd__clkinv_8 c622(
.A(net685),
.Y(out4)
);

sky130_fd_sc_hd__nor3_2 c623(
.A(net317),
.B(out19),
.C(net378),
.Y(net485)
);

sky130_fd_sc_hd__buf_16 c624(
.A(net687),
.X(net486)
);

sky130_fd_sc_hd__and3b_2 c625(
.A_N(in10),
.B(net114),
.C(net381),
.X(net487)
);

sky130_fd_sc_hd__clkbuf_8 c626(
.A(net687),
.X(net488)
);

sky130_fd_sc_hd__and3b_4 c627(
.A_N(net278),
.B(net44),
.C(net463),
.X(net489)
);

sky130_fd_sc_hd__sdfbbp_1 c628(
.D(net381),
.RESET_B(net480),
.SCD(net485),
.SCE(net457),
.SET_B(net44),
.CLK(clk),
.Q(net490)
);

sky130_fd_sc_hd__sedfxbp_2 c629(
.D(net44),
.DE(net489),
.SCD(out4),
.SCE(net485),
.CLK(clk),
.Q(net492),
.Q_N(net491)
);

sky130_fd_sc_hd__sedfxtp_1 c630(
.D(net4),
.DE(net485),
.SCD(net484),
.SCE(net463),
.CLK(clk),
.Q(net493)
);

sky130_fd_sc_hd__a2111o_1 c631(
.A1(net481),
.A2(net493),
.B1(net365),
.C1(net378),
.D1(net316),
.X(net494)
);

sky130_fd_sc_hd__dfbbn_2 c632(
.D(net476),
.RESET_B(net491),
.SET_B(net382),
.CLK_N(clk),
.Q(net495)
);

sky130_fd_sc_hd__dfbbp_1 c633(
.D(net483),
.RESET_B(net495),
.SET_B(net484),
.CLK(clk),
.Q(out17)
);

sky130_fd_sc_hd__nor3_2 c634(
.A(net241),
.B(net492),
.C(in43),
.Y(net496)
);

sky130_fd_sc_hd__nor3_2 c635(
.A(net424),
.B(net280),
.C(net44),
.Y(net497)
);

sky130_fd_sc_hd__mux4_1 c636(
.A0(net486),
.A1(net496),
.A2(out2),
.A3(net497),
.S0(net485),
.S1(net484),
.X(net498)
);

sky130_fd_sc_hd__sedfxtp_2 c637(
.D(net497),
.DE(net485),
.SCD(net278),
.SCE(net381),
.CLK(clk),
.Q(net499)
);

sky130_fd_sc_hd__buf_8 c660(
.A(net622),
.X(net500)
);

sky130_fd_sc_hd__and2_2 c661(
.A(net392),
.B(net403),
.X(net501)
);

sky130_fd_sc_hd__or2_2 c662(
.A(net405),
.B(in6),
.X(net502)
);

sky130_fd_sc_hd__dlygate4sd1_1 c663(
.A(net621),
.X(net503)
);

sky130_fd_sc_hd__nand2_2 c664(
.A(in10),
.B(net79),
.Y(net504)
);

sky130_fd_sc_hd__dfrtp_2 c665(
.D(net503),
.RESET_B(net201),
.CLK(clk),
.Q(net505)
);

sky130_fd_sc_hd__dfrtp_4 c666(
.D(net504),
.RESET_B(net201),
.CLK(clk),
.Q(net506)
);

sky130_fd_sc_hd__nand2b_1 c667(
.A_N(net303),
.B(net412),
.Y(net507)
);

sky130_fd_sc_hd__nor2b_4 c668(
.A(net413),
.B_N(net196),
.Y(net508)
);

sky130_fd_sc_hd__nand3_2 c669(
.A(net505),
.B(net413),
.C(net392),
.Y(net509)
);

sky130_fd_sc_hd__nand2_4 c670(
.A(net501),
.B(net405),
.Y(net510)
);

sky130_fd_sc_hd__dfsbp_1 c671(
.D(net201),
.SET_B(net292),
.CLK(clk),
.Q(net512),
.Q_N(net511)
);

sky130_fd_sc_hd__dfsbp_2 c672(
.D(net506),
.SET_B(net294),
.CLK(clk),
.Q(net514),
.Q_N(net513)
);

sky130_fd_sc_hd__or2_1 c673(
.A(in5),
.B(net505),
.X(net515)
);

sky130_fd_sc_hd__or2_2 c674(
.A(net403),
.B(net511),
.X(net516)
);

sky130_fd_sc_hd__or2b_4 c675(
.A(net514),
.B_N(net515),
.X(net517)
);

sky130_fd_sc_hd__dfstp_1 c676(
.D(net509),
.SET_B(net517),
.CLK(clk),
.Q(net518)
);

sky130_fd_sc_hd__and2b_4 c677(
.A_N(net507),
.B(net518),
.X(net519)
);

sky130_fd_sc_hd__and2_4 c678(
.A(net502),
.B(net505),
.X(net520)
);

sky130_fd_sc_hd__nand2b_1 c679(
.A_N(net518),
.B(net513),
.Y(net521)
);

sky130_fd_sc_hd__or2_4 c680(
.A(net521),
.B(net518),
.X(net522)
);

sky130_fd_sc_hd__sedfxtp_4 c681(
.D(net519),
.DE(net520),
.SCD(net508),
.SCE(net522),
.CLK(clk),
.Q(net523)
);

sky130_fd_sc_hd__nor3b_2 c682(
.A(net514),
.B(net431),
.C_N(net523),
.Y(net524)
);

sky130_fd_sc_hd__clkinv_1 c683(
.A(net626),
.Y(net525)
);

sky130_fd_sc_hd__nor2_1 c684(
.A(net427),
.B(net515),
.Y(net526)
);

sky130_fd_sc_hd__sdfxbp_1 c685(
.D(net503),
.SCD(out22),
.SCE(net216),
.CLK(clk),
.Q(net527)
);

sky130_fd_sc_hd__clkinv_16 c686(
.A(net625),
.Y(net528)
);

sky130_fd_sc_hd__inv_8 c687(
.Y(net529)
);

sky130_fd_sc_hd__and3_2 c688(
.A(net500),
.B(net516),
.C(net503),
.X(net530)
);

sky130_fd_sc_hd__nand3b_2 c689(
.A_N(net284),
.B(net510),
.C(net516),
.Y(net531)
);

sky130_fd_sc_hd__nand3_4 c690(
.A(net428),
.B(net512),
.C(net522),
.Y(net532)
);

sky130_fd_sc_hd__sdfxbp_2 c691(
.D(net532),
.SCD(net393),
.SCE(net528),
.CLK(clk),
.Q(net533)
);

sky130_fd_sc_hd__inv_6 c692(
.A(net649),
.Y(net534)
);

sky130_fd_sc_hd__sdfxtp_1 c693(
.D(net515),
.SCD(net294),
.SCE(net531),
.CLK(clk),
.Q(net535)
);

sky130_fd_sc_hd__nor3_1 c694(
.A(net534),
.B(net533),
.C(net284),
.Y(net536)
);

sky130_fd_sc_hd__nand2_4 c695(
.A(net535),
.B(net425),
.Y(net537)
);

sky130_fd_sc_hd__nor3_2 c696(
.A(net391),
.B(net535),
.C(net428),
.Y(net538)
);

sky130_fd_sc_hd__and2b_2 c697(
.A_N(net512),
.B(net500),
.X(net539)
);

sky130_fd_sc_hd__sdfxtp_2 c698(
.D(net531),
.SCD(in20),
.SCE(net196),
.CLK(clk),
.Q(net540)
);

sky130_fd_sc_hd__sdfxtp_4 c699(
.D(net294),
.SCD(net527),
.SCE(net427),
.CLK(clk),
.Q(net541)
);

sky130_fd_sc_hd__nor3_2 c700(
.A(net523),
.B(net540),
.C(net539),
.Y(net542)
);

sky130_fd_sc_hd__and3b_1 c701(
.A_N(net537),
.B(net539),
.C(net535),
.X(net543)
);

sky130_fd_sc_hd__dfbbn_1 c702(
.D(net538),
.RESET_B(net541),
.SET_B(net531),
.CLK_N(clk),
.Q(net545),
.Q_N(net544)
);

sky130_fd_sc_hd__mux4_1 c703(
.A0(in6),
.A1(net542),
.A2(net545),
.A3(net543),
.S0(net528),
.S1(net535),
.X(net546)
);

sky130_fd_sc_hd__dlygate4sd3_1 c704(
.A(net615),
.X(net547)
);

sky130_fd_sc_hd__nor3b_2 c705(
.A(net345),
.B(net524),
.C_N(net393),
.Y(net548)
);

sky130_fd_sc_hd__or3b_1 c706(
.A(net517),
.B(net539),
.C_N(net457),
.X(net549)
);

sky130_fd_sc_hd__nand2b_4 c707(
.A_N(net547),
.B(net121),
.Y(net550)
);

sky130_fd_sc_hd__dfbbn_2 c708(
.D(net301),
.RESET_B(net549),
.SET_B(net544),
.CLK_N(clk),
.Q(net552),
.Q_N(net551)
);

sky130_fd_sc_hd__and3b_1 c709(
.A_N(net425),
.B(net540),
.C(net547),
.X(net553)
);

sky130_fd_sc_hd__buf_16 c710(
.A(net616),
.X(net554)
);

sky130_fd_sc_hd__and3b_1 c711(
.A_N(net553),
.B(net550),
.C(net59),
.X(net555)
);

sky130_fd_sc_hd__nor3b_2 c712(
.A(net516),
.B(net517),
.C_N(net524),
.Y(net556)
);

sky130_fd_sc_hd__o2111a_1 c713(
.A1(net114),
.A2(net455),
.B1(net196),
.C1(net539),
.D1(net524),
.X(net557)
);

sky130_fd_sc_hd__sdfbbn_1 c714(
.D(net216),
.RESET_B(net555),
.SCD(net425),
.SCE(net549),
.SET_B(net198),
.CLK_N(clk),
.Q(net559),
.Q_N(net558)
);

sky130_fd_sc_hd__nor3_4 c715(
.A(net556),
.B(net393),
.C(net550),
.Y(net560)
);

sky130_fd_sc_hd__dfbbp_1 c716(
.D(net557),
.RESET_B(net549),
.SET_B(net216),
.CLK(clk),
.Q(net562),
.Q_N(net561)
);

sky130_fd_sc_hd__or4bb_1 c717(
.A(net520),
.B(net562),
.C_N(net453),
.D_N(net550),
.X(net563)
);

sky130_fd_sc_hd__nor3_2 c718(
.A(net559),
.B(in34),
.C(net524),
.Y(net564)
);

sky130_fd_sc_hd__or3_1 c719(
.A(net564),
.B(net524),
.C(net550),
.X(net565)
);

sky130_fd_sc_hd__sdfxbp_1 c720(
.D(net540),
.SCD(net453),
.SCE(net549),
.CLK(clk),
.Q(net567),
.Q_N(net566)
);

sky130_fd_sc_hd__mux4_4 c721(
.A0(net543),
.A1(net453),
.A2(net551),
.A3(net216),
.S0(net528),
.S1(net566),
.X(net568)
);

sky130_fd_sc_hd__nor3_2 c722(
.A(net425),
.B(net543),
.C(net672),
.Y(net569)
);

sky130_fd_sc_hd__or4bb_1 c723(
.A(net510),
.B(net550),
.C_N(net454),
.D_N(net569),
.X(net570)
);

sky130_fd_sc_hd__sdfxbp_2 c724(
.D(net567),
.SCD(net549),
.SCE(net558),
.CLK(clk),
.Q(net571)
);

sky130_fd_sc_hd__mux4_4 c725(
.A0(net536),
.A1(net565),
.A2(net292),
.A3(net561),
.S0(net549),
.S1(net569),
.X(net572)
);

sky130_fd_sc_hd__mux4_2 c726(
.A0(net198),
.A1(in59),
.A2(net393),
.A3(in5),
.S0(net528),
.S1(net554),
.X(net573)
);

sky130_fd_sc_hd__inv_6 c727(
.A(net686),
.Y(net574)
);

sky130_fd_sc_hd__inv_6 c728(
.A(net686),
.Y(net575)
);

sky130_fd_sc_hd__nand3b_4 c729(
.A_N(net196),
.B(net524),
.C(net85),
.Y(net576)
);

sky130_fd_sc_hd__sdfxtp_1 c730(
.D(net526),
.SCD(net570),
.SCE(in38),
.CLK(clk),
.Q(net577)
);

sky130_fd_sc_hd__mux4_1 c731(
.A0(net352),
.A1(net393),
.A2(in38),
.A3(net522),
.S0(net198),
.S1(net524),
.X(net578)
);

sky130_fd_sc_hd__or4bb_4 c732(
.A(net113),
.B(net545),
.C_N(net522),
.D_N(net198),
.X(net579)
);

sky130_fd_sc_hd__nand3_2 c733(
.A(net478),
.B(net548),
.C(net670),
.Y(net580)
);

sky130_fd_sc_hd__or4bb_4 c734(
.A(net262),
.B(net571),
.C_N(net352),
.D_N(net530),
.X(net581)
);

sky130_fd_sc_hd__sdfxtp_2 c735(
.D(net450),
.SCD(net459),
.SCE(net85),
.CLK(clk),
.Q(net582)
);

sky130_fd_sc_hd__mux4_2 c736(
.A0(net292),
.A1(net581),
.A2(net574),
.A3(net352),
.S0(net579),
.S1(net59),
.X(net583)
);

sky130_fd_sc_hd__sdfxtp_4 c737(
.D(net563),
.SCD(net569),
.SCE(net580),
.CLK(clk),
.Q(net584)
);

sky130_fd_sc_hd__nor3b_1 c738(
.A(net580),
.B(net578),
.C_N(net393),
.Y(net585)
);

sky130_fd_sc_hd__or3b_1 c739(
.A(net552),
.B(net585),
.C_N(net352),
.X(net586)
);

sky130_fd_sc_hd__a2111o_2 c740(
.A1(net85),
.A2(net575),
.B1(net580),
.C1(net585),
.D1(net123),
.X(net587)
);

sky130_fd_sc_hd__mux4_4 c741(
.A0(net554),
.A1(net584),
.A2(net586),
.A3(net292),
.S0(net198),
.S1(net352),
.X(net588)
);

sky130_fd_sc_hd__nand3b_4 c742(
.A_N(net479),
.B(net579),
.C(net576),
.Y(net589)
);

sky130_fd_sc_hd__dfbbn_1 c743(
.D(net522),
.RESET_B(net587),
.SET_B(net675),
.CLK_N(clk),
.Q(net590)
);

sky130_fd_sc_hd__and3b_1 c744(
.A_N(net263),
.B(net573),
.C(net589),
.X(net591)
);

sky130_fd_sc_hd__dfbbn_2 c745(
.D(net555),
.RESET_B(out0),
.SET_B(net676),
.CLK_N(clk),
.Q(net592)
);

sky130_fd_sc_hd__and3_1 c746(
.A(net590),
.B(net530),
.C(net592),
.X(net593)
);

sky130_fd_sc_hd__dfbbp_1 c747(
.D(net591),
.RESET_B(net593),
.SET_B(net368),
.CLK(clk),
.Q(net594)
);

sky130_fd_sc_hd__mux4_4 c748(
.A0(net560),
.A1(net548),
.A2(net499),
.A3(net85),
.S0(net589),
.S1(net436),
.X(net595)
);

sky130_fd_sc_hd__mux4_1 c749(
.A0(net453),
.A1(net435),
.A2(net121),
.A3(net589),
.S0(out22),
.S1(net674),
.X(net596)
);

sky130_fd_sc_hd__mux4_2 c750(
.A0(net596),
.A1(net382),
.A2(net482),
.A3(net589),
.S0(net387),
.S1(net673),
.X(net597)
);

sky130_fd_sc_hd__mux4_4 c751(
.A0(net494),
.A1(net378),
.A2(net582),
.A3(net560),
.S0(net85),
.S1(net589),
.X(net598)
);

sky130_fd_sc_hd__mux4_1 c752(
.A0(net457),
.A1(net589),
.A2(net301),
.A3(net387),
.S0(net677),
.S1(net679),
.X(net599)
);

sky130_fd_sc_hd__mux4_1 c753(
.A0(net577),
.A1(net387),
.A2(net599),
.A3(net59),
.S0(net85),
.S1(net671),
.X(net600)
);

sky130_fd_sc_hd__mux4_1 c754(
.A0(net477),
.A1(net436),
.A2(net594),
.A3(net59),
.S0(net589),
.S1(net680),
.X(net601)
);

sky130_fd_sc_hd__mux4_2 c755(
.A0(net490),
.A1(net488),
.A2(net599),
.A3(net589),
.S0(net678),
.S1(net681),
.X(net602)
);

sky130_fd_sc_hd__mux4_4 c756(
.A0(in53),
.A1(net487),
.A2(net589),
.A3(net680),
.S0(net681),
.S1(net682),
.X(net603)
);

sky130_fd_sc_hd__sdfrbp_1 merge757(
.D(net376),
.RESET_B(net271),
.Q(net377),
.SCE(out8),
.CLK(clk),
.Q_N(net604)
);

sky130_fd_sc_hd__sdfrbp_2 merge758(
.D(net247),
.RESET_B(net244),
.SCD(net110),
.SCE(net254),
.CLK(clk),
.Q(net607),
.Q_N(net606)
);

sky130_fd_sc_hd__sdfbbn_2 merge759(
.D(net268),
.RESET_B(net277),
.SCD(net260),
.SCE(net187),
.SET_B(net44),
.CLK_N(clk),
.Q(net609),
.Q_N(net608)
);

sky130_fd_sc_hd__sdfbbp_1 merge760(
.D(net150),
.RESET_B(net15),
.SCD(net29),
.SCE(out8),
.SET_B(net31),
.CLK(clk),
.Q(net611),
.Q_N(net610)
);

sky130_fd_sc_hd__sdfrtn_1 merge761(
.D(net217),
.RESET_B(net436),
.SCD(out14),
.SCE(net662),
.CLK_N(clk),
.Q(net612)
);

sky130_fd_sc_hd__sdfrtp_1 merge762(
.D(net308),
.RESET_B(net340),
.SCD(net358),
.SCE(net359),
.CLK(clk),
.Q(net613)
);

sky130_fd_sc_hd__mux4_1 merge763(
.A0(net88),
.A1(net197),
.A2(net211),
.A3(net218),
.S0(net214),
.S1(net219),
.X(net614)
);

sky130_fd_sc_hd__sdfbbn_1 merge764(
.D(net539),
.RESET_B(net319),
.SCD(net123),
.SCE(net520),
.SET_B(net216),
.CLK_N(clk),
.Q(net616),
.Q_N(net615)
);

sky130_fd_sc_hd__sdfrtp_2 merge765(
.D(net143),
.RESET_B(out1),
.SCD(net174),
.SCE(net173),
.CLK(clk),
.Q(net617)
);

sky130_fd_sc_hd__sdfrtp_4 merge766(
.D(net126),
.RESET_B(out46),
.SCD(net125),
.SCE(net2),
.CLK(clk),
.Q(net618)
);

sky130_fd_sc_hd__sdfbbn_2 merge767(
.D(net38),
.RESET_B(net36),
.Q(net40),
.SCE(net14),
.SET_B(net29),
.CLK_N(clk),
.Q_N(net619)
);

sky130_fd_sc_hd__sdfsbp_1 merge768(
.D(net294),
.SCD(net392),
.SCE(net412),
.SET_B(net201),
.CLK(clk),
.Q(net622),
.Q_N(net621)
);

sky130_fd_sc_hd__sdfsbp_2 merge769(
.D(net310),
.SCD(net287),
.SCE(net314),
.SET_B(net315),
.CLK(clk),
.Q(net624),
.Q_N(net623)
);

sky130_fd_sc_hd__sdfxbp_1 merge770(
.D(net79),
.SCD(net508),
.SCE(net198),
.CLK(clk),
.Q(net626),
.Q_N(net625)
);

sky130_fd_sc_hd__sdfbbp_1 merge771(
.D(net330),
.RESET_B(net302),
.SCD(in58),
.SCE(net332),
.SET_B(net338),
.CLK(clk),
.Q(net628),
.Q_N(net627)
);

sky130_fd_sc_hd__sdfstp_1 merge772(
.D(net359),
.SCD(net336),
.SCE(net264),
.SET_B(net465),
.CLK(clk),
.Q(net629)
);

sky130_fd_sc_hd__sdfbbn_1 merge773(
.D(net207),
.RESET_B(in58),
.SCD(net211),
.SCE(in49),
.SET_B(net226),
.CLK_N(clk),
.Q(net631),
.Q_N(net630)
);

sky130_fd_sc_hd__sdfstp_2 merge774(
.D(net395),
.SCD(net396),
.Q(net397),
.SET_B(net201),
.CLK(clk)
);

sky130_fd_sc_hd__sdfstp_4 merge775(
.D(net409),
.SCD(net216),
.SCE(net314),
.SET_B(net661),
.CLK(clk),
.Q(net633)
);

sky130_fd_sc_hd__mux4_4 merge776(
.A0(net463),
.A1(net301),
.A2(net382),
.A3(net298),
.S0(net390),
.S1(net457),
.X(net634)
);

sky130_fd_sc_hd__sedfxbp_1 merge777(
.D(net38),
.DE(out1),
.SCD(net41),
.SCE(net46),
.CLK(clk),
.Q(net636),
.Q_N(net635)
);

sky130_fd_sc_hd__mux4_2 merge778(
.A0(net393),
.A1(net546),
.A2(net563),
.A3(net528),
.S0(net368),
.S1(net522),
.X(net637)
);

sky130_fd_sc_hd__mux4_4 merge779(
.A0(net484),
.A1(net80),
.A2(in59),
.A3(net254),
.S0(net381),
.S1(out3),
.X(net638)
);

sky130_fd_sc_hd__sdfbbn_2 merge780(
.D(net43),
.RESET_B(out1),
.SCD(net126),
.SCE(in49),
.SET_B(in53),
.CLK_N(clk),
.Q(net640),
.Q_N(net639)
);

sky130_fd_sc_hd__mux4_1 merge781(
.A0(net219),
.A1(net372),
.A2(out7),
.A3(net177),
.S0(net173),
.S1(net172),
.X(net641)
);

sky130_fd_sc_hd__sedfxbp_2 merge782(
.D(net422),
.DE(net446),
.SCD(net93),
.SCE(net430),
.CLK(clk),
.Q(net643),
.Q_N(net642)
);

sky130_fd_sc_hd__sedfxtp_1 merge783(
.D(net293),
.DE(net291),
.SCD(net64),
.SCE(net310),
.CLK(clk),
.Q(net644)
);

sky130_fd_sc_hd__mux4_4 merge784(
.A0(net373),
.A1(net277),
.A2(net377),
.A3(net375),
.S0(net271),
.S1(net278),
.X(net645)
);

sky130_fd_sc_hd__sedfxtp_2 merge785(
.D(net448),
.DE(net216),
.SCD(net469),
.SCE(net470),
.CLK(clk),
.Q(net646)
);

sky130_fd_sc_hd__mux4_1 merge786(
.A0(net34),
.A1(in43),
.A2(net260),
.A3(in53),
.S0(net219),
.S1(in34),
.X(net647)
);

sky130_fd_sc_hd__sdfxbp_2 merge787(
.Q_N(net529),
.SCD(net319),
.SCE(net525),
.CLK(clk),
.Q(net649)
);

sky130_fd_sc_hd__mux4_4 merge788(
.A0(net221),
.A1(net240),
.A2(net242),
.A3(net237),
.S0(net238),
.S1(net235),
.X(net650)
);

sky130_fd_sc_hd__inv_1 merge789(
.A(net695),
.Y(net651)
);

sky130_fd_sc_hd__mux4_1 merge790(
.A0(net171),
.A1(net175),
.A2(out1),
.A3(net167),
.S0(net177),
.S1(net173),
.X(net652)
);

sky130_fd_sc_hd__sedfxtp_4 merge791(
.D(in20),
.DE(net201),
.SCD(net293),
.SCE(in3),
.CLK(clk),
.Q(net653)
);

sky130_fd_sc_hd__mux4_4 merge792(
.A0(net181),
.A1(net260),
.A2(net259),
.A3(net276),
.S0(net272),
.S1(out3),
.X(net654)
);

sky130_fd_sc_hd__sdfrbp_1 merge793(
.D(net249),
.RESET_B(net256),
.SCD(net332),
.SCE(net444),
.CLK(clk),
.Q(net656),
.Q_N(net655)
);

sky130_fd_sc_hd__dfxbp_1 s794(
.D(net163),
.CLK(clk),
.Q(out54),
.Q_N(net657)
);

sky130_fd_sc_hd__dfxbp_2 s795(
.D(net180),
.CLK(clk),
.Q(net658)
);

sky130_fd_sc_hd__dfxtp_1 s796(
.D(net202),
.CLK(clk),
.Q(out52)
);

sky130_fd_sc_hd__dfxtp_2 s797(
.D(net246),
.CLK(clk),
.Q(net659)
);

sky130_fd_sc_hd__dfxtp_4 s798(
.D(net281),
.CLK(clk),
.Q(out24)
);

sky130_fd_sc_hd__dlclkp_1 s799(
.GATE(net282),
.CLK(clk),
.GCLK(out34)
);

sky130_fd_sc_hd__dlclkp_2 s800(
.GATE(net305),
.CLK(clk),
.GCLK(net660)
);

sky130_fd_sc_hd__dlclkp_4 s801(
.GATE(net325),
.CLK(clk),
.GCLK(net661)
);

sky130_fd_sc_hd__dlxbn_1 s802(
.D(net327),
.GATE_N(clk),
.Q(net663),
.Q_N(net662)
);

sky130_fd_sc_hd__dlxbn_2 s803(
.D(net344),
.GATE_N(clk),
.Q(net665),
.Q_N(net664)
);

sky130_fd_sc_hd__dlxbp_1 s804(
.D(net347),
.GATE(clk),
.Q(net667),
.Q_N(net666)
);

sky130_fd_sc_hd__dlxtn_1 s805(
.D(net362),
.GATE_N(clk),
.Q(net668)
);

sky130_fd_sc_hd__dlxtn_2 s806(
.D(net458),
.GATE_N(clk),
.Q(net669)
);

sky130_fd_sc_hd__dlxtn_4 s807(
.D(net474),
.GATE_N(clk),
.Q(net670)
);

sky130_fd_sc_hd__dlxtp_1 s808(
.D(net498),
.GATE(clk),
.Q(net671)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s809(
.D(net568),
.SLEEP_B(clk),
.Q(net672)
);

sky130_fd_sc_hd__dfxbp_1 s810(
.D(net572),
.CLK(clk),
.Q(net674),
.Q_N(net673)
);

sky130_fd_sc_hd__dfxbp_2 s811(
.D(net583),
.CLK(clk),
.Q(net675)
);

sky130_fd_sc_hd__dfxtp_1 s812(
.D(net588),
.CLK(clk),
.Q(net676)
);

sky130_fd_sc_hd__dfxtp_2 s813(
.D(net595),
.CLK(clk),
.Q(net677)
);

sky130_fd_sc_hd__dfxtp_4 s814(
.D(net597),
.CLK(clk),
.Q(net678)
);

sky130_fd_sc_hd__dlclkp_1 s815(
.GATE(net598),
.CLK(clk),
.GCLK(net679)
);

sky130_fd_sc_hd__dlclkp_2 s816(
.GATE(net600),
.CLK(clk),
.GCLK(net680)
);

sky130_fd_sc_hd__dlclkp_4 s817(
.GATE(net601),
.CLK(clk),
.GCLK(net681)
);

sky130_fd_sc_hd__dlxbn_1 s818(
.D(net602),
.GATE_N(clk),
.Q(net682)
);

sky130_fd_sc_hd__dlxbn_2 s819(
.D(net603),
.GATE_N(clk)
);

sky130_fd_sc_hd__dlxbp_1 s820(
.D(net614),
.GATE(clk),
.Q(net684),
.Q_N(net683)
);

sky130_fd_sc_hd__dlxtn_1 s821(
.D(net634),
.GATE_N(clk),
.Q(net685)
);

sky130_fd_sc_hd__dlxtn_2 s822(
.D(net637),
.GATE_N(clk),
.Q(net686)
);

sky130_fd_sc_hd__dlxtn_4 s823(
.D(net638),
.GATE_N(clk),
.Q(net687)
);

sky130_fd_sc_hd__dlxtp_1 s824(
.D(net641),
.GATE(clk),
.Q(net688)
);

sky130_fd_sc_hd__lpflow_inputisolatch_1 s825(
.D(net645),
.SLEEP_B(clk),
.Q(net689)
);

sky130_fd_sc_hd__dfxbp_1 s826(
.D(net647),
.CLK(clk),
.Q(net691),
.Q_N(net690)
);

sky130_fd_sc_hd__dfxbp_2 s827(
.D(net650),
.CLK(clk),
.Q(net693),
.Q_N(net692)
);

sky130_fd_sc_hd__dfxtp_1 s828(
.D(net652),
.CLK(clk),
.Q(net694)
);

sky130_fd_sc_hd__dfxtp_2 s829(
.D(net654),
.CLK(clk),
.Q(net695)
);


endmodule
